`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  reg [34:0] PI_io_inputs;
  wire [0:0] PI_clock = clock;
  Sodor1StageTop UUT (
    .io_inputs(PI_io_inputs),
    .clock(PI_clock)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$formal$Sodor1Stage_formal.\sv:427$1_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:428$2_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:429$3_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:430$4_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:431$5_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:432$6_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:433$7_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:434$8_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:435$9_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:436$10_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:437$11_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:438$12_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:439$13_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:440$14_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:441$15_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:442$16_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:443$17_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:444$18_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:445$19_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:446$20_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:447$21_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:448$22_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:449$23_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:450$24_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:451$25_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:452$26_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:453$27_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:454$28_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:455$29_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:456$30_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:457$31_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:458$32_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:459$33_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:460$34_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:461$35_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:462$36_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:463$37_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:464$38_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:465$39_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:466$40_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:467$41_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:468$42_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:469$43_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:470$44_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:471$45_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:472$46_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:473$47_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:474$48_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:475$49_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:476$50_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:477$51_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:478$52_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:479$53_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:480$54_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:481$55_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:482$56_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:483$57_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:484$58_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:485$59_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:486$60_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:487$61_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:488$62_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:489$63_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:490$64_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:491$65_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:492$66_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:493$67_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:494$68_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:495$69_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:496$70_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:497$71_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:498$72_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:499$73_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:500$74_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:501$75_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:502$76_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:503$77_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:504$78_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:505$79_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:506$80_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:507$81_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:508$82_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:509$83_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:510$84_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:511$85_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:512$86_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:513$87_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:514$88_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:515$89_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:516$90_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:517$91_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:518$92_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:519$93_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:520$94_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:521$95_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:522$96_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:523$97_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:524$98_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:525$99_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:526$100_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:527$101_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:528$102_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:529$103_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:530$104_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:531$105_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:532$106_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:533$107_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:534$108_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:535$109_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:536$110_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:537$111_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:538$112_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:539$113_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:540$114_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:541$115_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:542$116_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:543$117_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:544$118_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:545$119_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:546$120_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:547$121_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:548$122_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:549$123_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:550$124_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:551$125_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:552$126_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:553$127_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:554$128_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:555$129_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:556$130_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:557$131_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:558$132_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:559$133_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:560$134_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:561$135_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:562$136_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:563$137_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:564$138_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:565$139_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:566$140_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:567$141_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:568$142_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:569$143_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:570$144_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:571$145_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:572$146_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:573$147_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:574$148_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:575$149_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:576$150_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:577$151_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:578$152_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:579$153_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:580$154_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:581$155_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:582$156_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:583$157_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:584$158_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:585$159_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:586$160_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:587$161_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:588$162_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:589$163_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:590$164_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:591$165_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:592$166_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:593$167_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:594$168_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:595$169_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:596$170_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:597$171_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:598$172_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:599$173_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:600$174_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:601$175_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:602$176_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:603$177_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:604$178_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:605$179_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:606$180_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:607$181_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:608$182_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:609$183_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:610$184_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:611$185_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:612$186_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:613$187_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:614$188_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:615$189_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:616$190_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:617$191_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:618$192_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:619$193_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:620$194_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:621$195_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:622$196_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:623$197_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:624$198_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:625$199_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:626$200_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:627$201_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:628$202_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:629$203_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:630$204_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:631$205_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:632$206_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:633$207_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:634$208_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:635$209_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:636$210_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:637$211_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:638$212_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:639$213_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:640$214_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:641$215_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:642$216_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:643$217_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:644$218_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:645$219_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:646$220_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:647$221_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:648$222_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:649$223_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:650$224_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:651$225_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:652$226_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:653$227_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:654$228_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:655$229_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:656$230_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:657$231_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:658$232_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:659$233_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:660$234_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:661$235_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:662$236_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:663$237_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:664$238_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:665$239_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:666$240_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:667$241_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:668$242_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:669$243_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:670$244_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:671$245_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:672$246_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:673$247_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:674$248_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:675$249_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:676$250_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:677$251_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:678$252_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:679$253_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:680$254_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:681$255_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:682$256_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:683$257_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:684$258_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:685$259_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:686$260_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:687$261_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:688$262_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:689$263_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:690$264_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:691$265_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:692$266_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:693$267_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:694$268_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:695$269_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:696$270_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:697$271_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:698$272_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:699$273_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:700$274_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:701$275_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:702$276_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:703$277_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:704$278_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:705$279_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:706$280_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:707$281_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:708$282_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:709$283_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:710$284_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:711$285_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:712$286_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:713$287_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:714$288_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:715$289_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:716$290_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:717$291_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:718$292_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:719$293_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:720$294_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:721$295_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:722$296_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:723$297_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:724$298_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:725$299_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:726$300_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:727$301_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:728$302_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:729$303_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:730$304_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:731$305_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:732$306_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:733$307_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:734$308_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:735$309_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:736$310_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:737$311_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:738$312_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:739$313_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:740$314_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:741$315_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:742$316_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:743$317_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:744$318_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:745$319_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:746$320_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:747$321_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:748$322_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:749$323_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:750$324_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:751$325_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:752$326_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:753$327_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:754$328_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:755$329_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:756$330_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:757$331_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:758$332_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:759$333_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:760$334_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:761$335_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:762$336_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:763$337_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:764$338_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:765$339_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:766$340_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:767$341_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:768$342_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:769$343_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:770$344_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:771$345_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:772$346_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:773$347_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:774$348_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:775$349_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:776$350_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:777$351_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:778$352_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:779$353_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:780$354_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:781$355_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:782$356_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:783$357_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:784$358_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:785$359_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:786$360_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:787$361_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:788$362_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:789$363_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:790$364_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:791$365_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:792$366_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:793$367_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:794$368_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:795$369_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:796$370_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:797$371_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:798$372_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:799$373_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:800$374_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:801$375_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:802$376_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:803$377_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:804$378_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:805$379_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:806$380_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:807$381_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:808$382_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:809$383_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:810$384_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:811$385_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:812$386_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:813$387_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:814$388_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:815$389_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:816$390_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:817$391_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:818$392_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:819$393_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:820$394_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:821$395_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:822$396_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:823$397_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:824$398_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:825$399_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:826$400_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:827$401_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:828$402_CHECK  = 1'b0;
    // UUT.$formal$Sodor1Stage_formal.\sv:836$403_EN  = 1'b0;
    UUT.bb.core.d.csr._T_176 = 6'b111111;
    UUT.bb.core.d.csr._T_180 = 58'b0000000000000000000000000000000011111111111111111111111111;
    UUT.bb.core.d.csr._T_188 = 6'b111111;
    UUT.bb.core.d.csr._T_192 = 58'b0000000000000000000000000000000011111111111111111111111111;
    UUT.bb.core.d.csr._T_200 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_203 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_206 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_209 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_212 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_215 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_218 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_221 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_224 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_227 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_230 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_233 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_236 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_239 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_242 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_245 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_248 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_251 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_254 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_257 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_260 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_263 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_266 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_269 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_272 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_275 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_278 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_281 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_284 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_287 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_290 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr._T_293 = 40'b0000000011111111111111111111111111111111;
    UUT.bb.core.d.csr.reg_dcsr_ebreakm = 1'b1;
    UUT.bb.core.d.csr.reg_dcsr_step = 1'b1;
    UUT.bb.core.d.csr.reg_dpc = 32'b11111111111111111111111111111111;
    UUT.bb.core.d.csr.reg_dscratch = 32'b11111111111111111111111111111111;
    UUT.bb.core.d.csr.reg_mcause = 32'b11111111111111111111111111111111;
    UUT.bb.core.d.csr.reg_medeleg = 32'b11111111111111111111111111111111;
    UUT.bb.core.d.csr.reg_mepc = 32'b11111111111111111111111111111111;
    UUT.bb.core.d.csr.reg_mie_msip = 1'b1;
    UUT.bb.core.d.csr.reg_mie_mtip = 1'b1;
    UUT.bb.core.d.csr.reg_mip_msip = 1'b1;
    UUT.bb.core.d.csr.reg_mip_mtip = 1'b1;
    UUT.bb.core.d.csr.reg_mscratch = 32'b11111111111111111111111111111111;
    UUT.bb.core.d.csr.reg_mstatus_mie = 1'b1;
    UUT.bb.core.d.csr.reg_mstatus_mpie = 1'b1;
    UUT.bb.core.d.csr.reg_mtval = 32'b11111111111111111111111111111111;
    UUT.bb.core.d.mem_sparse.addresses_0_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_0_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_10_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_10_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_11_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_11_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_12_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_12_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_13_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_13_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_14_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_14_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_15_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_15_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_16_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_16_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_17_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_17_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_18_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_18_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_19_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_19_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_1_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_1_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_20_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_20_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_21_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_21_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_22_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_22_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_23_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_23_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_24_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_24_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_25_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_25_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_26_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_26_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_27_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_27_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_28_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_28_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_29_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_29_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_2_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_2_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_30_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_30_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_31_bits = 5'b10000;
    UUT.bb.core.d.mem_sparse.addresses_31_valid = 1'b1;
    UUT.bb.core.d.mem_sparse.addresses_3_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_3_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_4_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_4_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_5_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_5_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_6_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_6_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_7_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_7_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_8_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_8_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.addresses_9_bits = 5'b00000;
    UUT.bb.core.d.mem_sparse.addresses_9_valid = 1'b0;
    UUT.bb.core.d.mem_sparse.nextAddr = 6'b100000;
    UUT.bb.core.d.pc_reg = 32'b11111111111111111111111111110111;
    UUT.bb.memory.async_data.mem_sparse.addresses_0_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_10_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_11_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_12_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_13_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_14_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_15_bits = 21'b000000000000000000000;
    UUT.bb.memory.async_data.mem_sparse.addresses_16_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_17_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_18_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_19_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_1_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_20_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_21_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_22_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_23_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_24_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_25_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_26_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_27_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_28_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_29_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_2_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_30_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_31_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_3_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_4_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_5_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_6_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_7_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_8_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_9_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.nextAddr = 6'b111110;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_0_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_10_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_11_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_12_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_13_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_14_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_15_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_16_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_17_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_18_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_19_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_1_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_20_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_21_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_22_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_23_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_24_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_25_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_26_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_27_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_28_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_29_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_2_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_30_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_31_bits = 21'b000000000000000000000;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_3_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_4_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_5_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_6_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_7_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_8_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_9_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.nextAddr = 6'b111110;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_0_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_10_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_11_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_12_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_13_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_14_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_15_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_16_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_17_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_18_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_19_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_1_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_20_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_21_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_22_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_23_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_24_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_25_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_26_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_27_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_28_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_29_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_2_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_30_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_31_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_3_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_4_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_5_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_6_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_7_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_8_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_9_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.nextAddr = 6'b111110;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_0_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_10_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_11_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_12_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_13_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_14_bits = 21'b000000000000000000000;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_15_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_16_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_17_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_18_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_19_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_1_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_20_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_21_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_22_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_23_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_24_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_25_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_26_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_27_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_28_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_29_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_2_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_30_bits = 21'b000000000000000000000;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_31_bits = 21'b000000000000000000011;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_3_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_4_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_5_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_6_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_7_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_8_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_9_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.nextAddr = 6'b111110;
    UUT.is_meta_reset_phase = 1'b1;
    UUT.is_reset_phase = 1'b0;
    UUT.bb.core.d.mem_sparse.mem[5'b11111] = 32'b00000000011111111111111011111111;
    UUT.bb.core.d.mem_sparse.mem[5'b00000] = 32'b00000000000000000000000000000000;
    UUT.bb.memory.async_data.mem_sparse.mem[5'b01111] = 8'b00000000;
    UUT.bb.memory.async_data.mem_sparse.mem[5'b00000] = 8'b11111111;
    UUT.bb.memory.async_data.mem_sparse.mem[5'b11111] = 8'b11111111;
    UUT.bb.memory.async_data.mem_sparse_0.mem[5'b11111] = 8'b11111111;
    UUT.bb.memory.async_data.mem_sparse_0.mem[5'b00000] = 8'b11111111;
    UUT.bb.memory.async_data.mem_sparse_1.mem[5'b11111] = 8'b11111111;
    UUT.bb.memory.async_data.mem_sparse_1.mem[5'b00000] = 8'b11111111;
    UUT.bb.memory.async_data.mem_sparse_2.mem[5'b11111] = 8'b11111111;
    UUT.bb.memory.async_data.mem_sparse_2.mem[5'b00000] = 8'b11111111;

    // state 0
    PI_io_inputs = 35'b10001111000010000011000000010011010;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_io_inputs <= 35'b00000000000100000000000000010111010;
    end

    // state 2
    if (cycle == 1) begin
      PI_io_inputs <= 35'b10110000110000001000100000001111010;
    end

    // state 3
    if (cycle == 2) begin
      PI_io_inputs <= 35'b10000000000111110010111110010011010;
    end

    genclock <= cycle < 3;
    cycle <= cycle + 1;
  end
endmodule
