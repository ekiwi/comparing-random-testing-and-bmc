`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  wire [0:0] PI_clock = clock;
  TileAndMemTop UUT (
    .clock(PI_clock)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    UUT._resetCount = 1'b0;
    UUT.addr = 32'b00000000000000000000000000000000;
    UUT.dut.arb.state = 3'b000;
    UUT.dut.core.dpath.csr.IE = 1'b0;
    UUT.dut.core.dpath.csr.IE1 = 1'b0;
    UUT.dut.core.dpath.csr.MSIE = 1'b0;
    UUT.dut.core.dpath.csr.MSIP = 1'b0;
    UUT.dut.core.dpath.csr.MTIE = 1'b0;
    UUT.dut.core.dpath.csr.MTIP = 1'b0;
    UUT.dut.core.dpath.csr.PRV = 2'b00;
    UUT.dut.core.dpath.csr.PRV1 = 2'b00;
    UUT.dut.core.dpath.csr.cycle = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.cycleh = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.instret = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.instreth = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.mbadaddr = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.mcause = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.mepc = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.mfromhost = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.mscratch = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.mtimecmp = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.mtohost = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.time_ = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr.timeh = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.csr_cmd = 3'b000;
    UUT.dut.core.dpath.csr_in = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.ew_alu = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.ew_inst = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.ew_pc = 33'b000000000000000000000000000000000;
    UUT.dut.core.dpath.fe_inst = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.fe_pc = 33'b000000000000000000000000000000000;
    UUT.dut.core.dpath.illegal = 1'b0;
    UUT.dut.core.dpath.ld_type = 3'b000;
    UUT.dut.core.dpath.pc = 33'b000000000000000000000000000000000;
    UUT.dut.core.dpath.pc_check = 1'b0;
    UUT.dut.core.dpath.st_type = 2'b00;
    UUT.dut.core.dpath.started = 1'b0;
    UUT.dut.core.dpath.wb_en = 1'b0;
    UUT.dut.core.dpath.wb_sel = 2'b00;
    UUT.dut.dcache.addr_reg = 32'b00000000000000000000000000000000;
    UUT.dut.dcache.cpu_data = 32'b00000000000000000000000000000000;
    UUT.dut.dcache.cpu_mask = 4'b0000;
    UUT.dut.dcache.d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.dcache.dataMem_3_3_rdata_MPORT_3_addr_pipe_0 = 8'b00000000;
    UUT.dut.dcache.is_alloc_reg = 1'b0;
    UUT.dut.dcache.rdata_buf = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.dcache.read_count = 1'b0;
    UUT.dut.dcache.refill_buf_0 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.dcache.refill_buf_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.dcache.ren_reg = 1'b0;
    UUT.dut.dcache.state = 3'b000;
    UUT.dut.dcache.v = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.dcache.write_count = 1'b0;
    UUT.dut.icache.addr_reg = 32'b00000000000000000000000000000000;
    UUT.dut.icache.d = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.icache.dataMem_3_3_rdata_MPORT_3_addr_pipe_0 = 8'b00000000;
    UUT.dut.icache.is_alloc_reg = 1'b0;
    UUT.dut.icache.rdata_buf = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.icache.read_count = 1'b0;
    UUT.dut.icache.refill_buf_0 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.icache.refill_buf_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.dut.icache.ren_reg = 1'b0;
    UUT.dut.icache.state = 3'b000;
    UUT.dut.icache.v = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.off = 8'b00000000;
    UUT.state = 2'b00;
    // UUT.tracker.$formal$SignalTracker.\sv:10001$3331_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10004$3332_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10007$3333_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1001$331_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10010$3334_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10013$3335_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10016$3336_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10019$3337_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10022$3338_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10025$3339_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10028$3340_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10031$3341_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10034$3342_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10037$3343_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1004$332_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10040$3344_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10043$3345_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10046$3346_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10049$3347_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10052$3348_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10055$3349_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10058$3350_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10061$3351_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10064$3352_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10067$3353_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1007$333_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10070$3354_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10073$3355_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10076$3356_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10079$3357_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10082$3358_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10085$3359_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10088$3360_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10091$3361_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10094$3362_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10097$3363_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1010$334_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10100$3364_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10103$3365_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10106$3366_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10109$3367_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10112$3368_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10115$3369_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10118$3370_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10121$3371_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10124$3372_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10127$3373_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1013$335_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10130$3374_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10133$3375_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10136$3376_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10139$3377_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10142$3378_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10145$3379_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10148$3380_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10151$3381_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10154$3382_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10157$3383_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1016$336_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10160$3384_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10163$3385_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10166$3386_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10169$3387_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10172$3388_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10175$3389_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10178$3390_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10181$3391_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10184$3392_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10187$3393_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1019$337_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10190$3394_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10193$3395_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10196$3396_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10199$3397_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10202$3398_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10205$3399_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10208$3400_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10211$3401_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10214$3402_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10217$3403_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1022$338_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10220$3404_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10223$3405_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10226$3406_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10229$3407_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10232$3408_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10235$3409_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10238$3410_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10241$3411_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10244$3412_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10247$3413_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1025$339_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10250$3414_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10253$3415_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10256$3416_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10259$3417_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10262$3418_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10265$3419_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10268$3420_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10271$3421_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10274$3422_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10277$3423_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1028$340_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10280$3424_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10283$3425_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10286$3426_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10289$3427_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10292$3428_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10295$3429_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10298$3430_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10301$3431_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10304$3432_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10307$3433_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1031$341_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10310$3434_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10313$3435_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10316$3436_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10319$3437_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10322$3438_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10325$3439_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10328$3440_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10331$3441_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10334$3442_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10337$3443_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1034$342_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10340$3444_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10343$3445_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10346$3446_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10349$3447_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10352$3448_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10355$3449_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10358$3450_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10361$3451_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10364$3452_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10367$3453_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1037$343_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10370$3454_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10373$3455_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10376$3456_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10379$3457_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10382$3458_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10385$3459_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10388$3460_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10391$3461_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10394$3462_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10397$3463_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1040$344_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10400$3464_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10403$3465_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10406$3466_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10409$3467_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10412$3468_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10415$3469_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10418$3470_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10421$3471_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10424$3472_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10427$3473_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1043$345_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10430$3474_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10433$3475_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10436$3476_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10439$3477_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10442$3478_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10445$3479_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10448$3480_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10451$3481_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10454$3482_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10457$3483_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1046$346_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10460$3484_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10463$3485_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10466$3486_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10469$3487_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10472$3488_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10475$3489_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10478$3490_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10481$3491_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10484$3492_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10487$3493_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1049$347_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10490$3494_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10493$3495_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10496$3496_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10499$3497_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10502$3498_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10505$3499_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10508$3500_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10511$3501_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10514$3502_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10517$3503_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1052$348_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10520$3504_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10523$3505_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10526$3506_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10529$3507_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10532$3508_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10535$3509_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10538$3510_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10541$3511_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10544$3512_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10547$3513_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1055$349_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10550$3514_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10553$3515_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10556$3516_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10559$3517_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10562$3518_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10565$3519_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10568$3520_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10571$3521_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10574$3522_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10577$3523_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1058$350_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10580$3524_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10583$3525_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10586$3526_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10589$3527_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10592$3528_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10595$3529_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10598$3530_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10601$3531_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10604$3532_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10607$3533_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1061$351_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10610$3534_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10613$3535_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10616$3536_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10619$3537_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10622$3538_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10625$3539_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10628$3540_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10631$3541_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10634$3542_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10637$3543_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1064$352_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10640$3544_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10643$3545_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10646$3546_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10649$3547_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10652$3548_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10655$3549_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10658$3550_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10661$3551_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10664$3552_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10667$3553_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1067$353_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10670$3554_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10673$3555_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10676$3556_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10679$3557_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10682$3558_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10685$3559_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10688$3560_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10691$3561_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10694$3562_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10697$3563_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1070$354_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10700$3564_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10703$3565_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10706$3566_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10709$3567_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10712$3568_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10715$3569_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10718$3570_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10721$3571_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10724$3572_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10727$3573_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1073$355_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10730$3574_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10733$3575_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10736$3576_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10739$3577_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10742$3578_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10745$3579_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10748$3580_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10751$3581_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10754$3582_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10757$3583_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1076$356_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10760$3584_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10763$3585_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10766$3586_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10769$3587_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10772$3588_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10775$3589_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10778$3590_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10781$3591_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10784$3592_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10787$3593_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1079$357_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10790$3594_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10793$3595_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10796$3596_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10799$3597_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10802$3598_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10805$3599_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10808$3600_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10811$3601_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10814$3602_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10817$3603_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1082$358_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10820$3604_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10823$3605_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10826$3606_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10829$3607_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10832$3608_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10835$3609_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10838$3610_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10841$3611_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10844$3612_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10847$3613_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1085$359_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10850$3614_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10853$3615_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10856$3616_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10859$3617_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10862$3618_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10865$3619_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10868$3620_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10871$3621_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10874$3622_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10877$3623_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1088$360_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10880$3624_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10883$3625_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10886$3626_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10889$3627_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10892$3628_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10895$3629_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10898$3630_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10901$3631_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10904$3632_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10907$3633_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1091$361_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10910$3634_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10913$3635_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10916$3636_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10919$3637_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10922$3638_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10925$3639_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10928$3640_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10931$3641_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10934$3642_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10937$3643_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1094$362_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10940$3644_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10943$3645_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10946$3646_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10949$3647_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10952$3648_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10955$3649_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10958$3650_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10961$3651_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10964$3652_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10967$3653_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1097$363_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10970$3654_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10973$3655_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10976$3656_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10979$3657_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10982$3658_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10985$3659_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10988$3660_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10991$3661_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10994$3662_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:10997$3663_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1100$364_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11000$3664_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11003$3665_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11006$3666_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11009$3667_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11012$3668_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11015$3669_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11018$3670_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11021$3671_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11024$3672_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11027$3673_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1103$365_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11030$3674_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11033$3675_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11036$3676_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11039$3677_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11042$3678_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11045$3679_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11048$3680_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11051$3681_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11054$3682_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11057$3683_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1106$366_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11060$3684_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11063$3685_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11066$3686_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11069$3687_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11072$3688_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11075$3689_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11078$3690_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11081$3691_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11084$3692_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11087$3693_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1109$367_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11090$3694_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11093$3695_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11096$3696_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11099$3697_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11102$3698_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11105$3699_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11108$3700_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11111$3701_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11114$3702_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11117$3703_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1112$368_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11120$3704_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11123$3705_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11126$3706_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11129$3707_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11132$3708_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11135$3709_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11138$3710_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11141$3711_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11144$3712_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11147$3713_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1115$369_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11150$3714_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11153$3715_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11156$3716_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11159$3717_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11162$3718_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11165$3719_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11168$3720_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11171$3721_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11174$3722_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11177$3723_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1118$370_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11180$3724_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11183$3725_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11186$3726_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11189$3727_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11192$3728_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11195$3729_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11198$3730_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11201$3731_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11204$3732_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11207$3733_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1121$371_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11210$3734_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11213$3735_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11216$3736_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11219$3737_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11222$3738_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11225$3739_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11228$3740_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11231$3741_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11234$3742_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11237$3743_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1124$372_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11240$3744_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11243$3745_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11246$3746_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11249$3747_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11252$3748_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11255$3749_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11258$3750_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11261$3751_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11264$3752_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11267$3753_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1127$373_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11270$3754_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11273$3755_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11276$3756_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11279$3757_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11282$3758_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11285$3759_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11288$3760_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11291$3761_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11294$3762_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11297$3763_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1130$374_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11300$3764_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11303$3765_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11306$3766_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11309$3767_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11312$3768_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11315$3769_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11318$3770_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11321$3771_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11324$3772_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11327$3773_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1133$375_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11330$3774_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11333$3775_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11336$3776_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11339$3777_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11342$3778_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11345$3779_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11348$3780_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11351$3781_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11354$3782_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11357$3783_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1136$376_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11360$3784_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11363$3785_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11366$3786_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11369$3787_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11372$3788_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11375$3789_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11378$3790_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11381$3791_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11384$3792_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11387$3793_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1139$377_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11390$3794_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11393$3795_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11396$3796_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11399$3797_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11402$3798_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11405$3799_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11408$3800_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11411$3801_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11414$3802_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11417$3803_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1142$378_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11420$3804_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11423$3805_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11426$3806_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11429$3807_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11432$3808_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11435$3809_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11438$3810_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11441$3811_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11444$3812_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11447$3813_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1145$379_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11450$3814_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11453$3815_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11456$3816_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11459$3817_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11462$3818_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11465$3819_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11468$3820_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11471$3821_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11474$3822_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11477$3823_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1148$380_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11480$3824_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11483$3825_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11486$3826_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11489$3827_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11492$3828_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11495$3829_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11498$3830_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11501$3831_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11504$3832_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11507$3833_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1151$381_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11510$3834_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11513$3835_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11516$3836_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11519$3837_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11522$3838_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11525$3839_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11528$3840_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11531$3841_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11534$3842_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11537$3843_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1154$382_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11540$3844_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11543$3845_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11546$3846_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11549$3847_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11552$3848_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11555$3849_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11558$3850_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11561$3851_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11564$3852_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11567$3853_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1157$383_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11570$3854_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11573$3855_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11576$3856_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11579$3857_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11582$3858_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11585$3859_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11588$3860_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11591$3861_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11594$3862_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11597$3863_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1160$384_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11600$3864_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11603$3865_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11606$3866_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11609$3867_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11612$3868_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11615$3869_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11618$3870_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11621$3871_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11624$3872_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11627$3873_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1163$385_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11630$3874_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11633$3875_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11636$3876_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11639$3877_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11642$3878_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11645$3879_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11648$3880_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11651$3881_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11654$3882_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11657$3883_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1166$386_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11660$3884_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11663$3885_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11666$3886_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11669$3887_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11672$3888_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11675$3889_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11678$3890_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11681$3891_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11684$3892_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11687$3893_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1169$387_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11690$3894_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11693$3895_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11696$3896_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11699$3897_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11702$3898_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11705$3899_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11708$3900_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11711$3901_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11714$3902_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11717$3903_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1172$388_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11720$3904_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11723$3905_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11726$3906_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11729$3907_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11732$3908_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11735$3909_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11738$3910_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11741$3911_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11744$3912_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11747$3913_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1175$389_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11750$3914_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11753$3915_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11756$3916_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11759$3917_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11762$3918_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11765$3919_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11768$3920_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11771$3921_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11774$3922_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11777$3923_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1178$390_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11780$3924_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11783$3925_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11786$3926_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11789$3927_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11792$3928_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11795$3929_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11798$3930_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11801$3931_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11804$3932_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11807$3933_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1181$391_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11810$3934_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11813$3935_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11816$3936_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11819$3937_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11822$3938_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11825$3939_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11828$3940_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11831$3941_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11834$3942_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11837$3943_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1184$392_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11840$3944_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11843$3945_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11846$3946_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11849$3947_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11852$3948_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11855$3949_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11858$3950_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11861$3951_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11864$3952_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11867$3953_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1187$393_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11870$3954_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11873$3955_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11876$3956_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11879$3957_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11882$3958_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11885$3959_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11888$3960_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11891$3961_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11894$3962_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11897$3963_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1190$394_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11900$3964_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11903$3965_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11906$3966_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11909$3967_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11912$3968_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11915$3969_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11918$3970_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11921$3971_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11924$3972_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11927$3973_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1193$395_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11930$3974_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11933$3975_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11936$3976_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11939$3977_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11942$3978_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11945$3979_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11948$3980_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11951$3981_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11954$3982_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11957$3983_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1196$396_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11960$3984_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11963$3985_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11966$3986_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11969$3987_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11972$3988_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11975$3989_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11978$3990_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11981$3991_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11984$3992_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11987$3993_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1199$397_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11990$3994_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11993$3995_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11996$3996_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:11999$3997_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12002$3998_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12005$3999_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12008$4000_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12011$4001_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12014$4002_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12017$4003_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1202$398_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12020$4004_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12023$4005_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12026$4006_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12029$4007_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12032$4008_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12035$4009_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12038$4010_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12041$4011_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12044$4012_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12047$4013_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1205$399_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12050$4014_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12053$4015_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12056$4016_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12059$4017_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12062$4018_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12065$4019_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12068$4020_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12071$4021_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12074$4022_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12077$4023_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1208$400_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12080$4024_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12083$4025_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12086$4026_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12089$4027_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12092$4028_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12095$4029_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12098$4030_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12101$4031_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12104$4032_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12107$4033_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1211$401_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12110$4034_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12113$4035_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12116$4036_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12119$4037_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12122$4038_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12125$4039_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12128$4040_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12131$4041_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12134$4042_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12137$4043_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1214$402_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12140$4044_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12143$4045_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12146$4046_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12149$4047_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12152$4048_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12155$4049_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12158$4050_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12161$4051_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12164$4052_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12167$4053_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1217$403_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12170$4054_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12173$4055_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12176$4056_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12179$4057_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12182$4058_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12185$4059_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12188$4060_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12191$4061_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12194$4062_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12197$4063_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1220$404_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12200$4064_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12203$4065_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12206$4066_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12209$4067_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12212$4068_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12215$4069_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12218$4070_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12221$4071_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12224$4072_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12227$4073_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1223$405_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12230$4074_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12233$4075_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12236$4076_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12239$4077_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12242$4078_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12245$4079_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12248$4080_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12251$4081_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12254$4082_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12257$4083_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1226$406_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12260$4084_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12263$4085_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12266$4086_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12269$4087_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12272$4088_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12275$4089_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12278$4090_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12281$4091_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12284$4092_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12287$4093_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1229$407_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12290$4094_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12293$4095_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12296$4096_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12299$4097_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12302$4098_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12305$4099_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12308$4100_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12311$4101_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12314$4102_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12317$4103_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1232$408_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12320$4104_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12323$4105_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12326$4106_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12329$4107_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12332$4108_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12335$4109_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12338$4110_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12341$4111_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12344$4112_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12347$4113_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1235$409_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12350$4114_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12353$4115_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12356$4116_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12359$4117_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12362$4118_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12365$4119_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12368$4120_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12371$4121_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12374$4122_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12377$4123_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1238$410_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12380$4124_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12383$4125_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12386$4126_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12389$4127_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12392$4128_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12395$4129_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12398$4130_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12401$4131_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12404$4132_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12407$4133_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1241$411_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12410$4134_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12413$4135_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12416$4136_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12419$4137_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12422$4138_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12425$4139_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12428$4140_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12431$4141_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12434$4142_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12437$4143_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1244$412_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12440$4144_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12443$4145_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12446$4146_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12449$4147_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12452$4148_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12455$4149_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12458$4150_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12461$4151_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12464$4152_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12467$4153_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1247$413_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12470$4154_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12473$4155_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12476$4156_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12479$4157_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12482$4158_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12485$4159_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12488$4160_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12491$4161_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12494$4162_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12497$4163_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1250$414_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12500$4164_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12503$4165_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12506$4166_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12509$4167_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12512$4168_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12515$4169_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12518$4170_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12521$4171_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12524$4172_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12527$4173_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1253$415_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12530$4174_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12533$4175_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12536$4176_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12539$4177_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12542$4178_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12545$4179_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12548$4180_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12551$4181_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12554$4182_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12557$4183_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1256$416_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12560$4184_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12563$4185_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12566$4186_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12569$4187_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12572$4188_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12575$4189_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12578$4190_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12581$4191_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12584$4192_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12587$4193_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1259$417_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12590$4194_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12593$4195_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12596$4196_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12599$4197_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12602$4198_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12605$4199_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12608$4200_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12611$4201_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12614$4202_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12617$4203_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1262$418_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12620$4204_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12623$4205_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12626$4206_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12629$4207_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12632$4208_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12635$4209_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12638$4210_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12641$4211_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12644$4212_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12647$4213_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1265$419_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12650$4214_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12653$4215_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12656$4216_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12659$4217_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12662$4218_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12665$4219_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12668$4220_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12671$4221_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12674$4222_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12677$4223_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1268$420_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12680$4224_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12683$4225_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12686$4226_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12689$4227_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12692$4228_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12695$4229_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12698$4230_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12701$4231_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12704$4232_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12707$4233_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1271$421_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12710$4234_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12713$4235_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12716$4236_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12719$4237_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12722$4238_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12725$4239_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12728$4240_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12731$4241_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12734$4242_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12737$4243_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1274$422_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12740$4244_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12743$4245_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12746$4246_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12749$4247_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12752$4248_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12755$4249_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12758$4250_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12761$4251_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12764$4252_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12767$4253_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1277$423_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12770$4254_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12773$4255_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12776$4256_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12779$4257_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12782$4258_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12785$4259_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12788$4260_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12791$4261_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12794$4262_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12797$4263_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1280$424_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12800$4264_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12803$4265_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12806$4266_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12809$4267_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12812$4268_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12815$4269_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12818$4270_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12821$4271_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12824$4272_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12827$4273_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1283$425_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12830$4274_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12833$4275_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12836$4276_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12839$4277_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12842$4278_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12845$4279_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12848$4280_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12851$4281_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12854$4282_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12857$4283_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1286$426_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12860$4284_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12863$4285_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12866$4286_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12869$4287_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12872$4288_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12875$4289_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12878$4290_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12881$4291_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12884$4292_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12887$4293_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1289$427_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12890$4294_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12893$4295_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12896$4296_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12899$4297_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12902$4298_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12905$4299_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12908$4300_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12911$4301_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12914$4302_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12917$4303_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1292$428_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12920$4304_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12923$4305_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12926$4306_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12929$4307_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12932$4308_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12935$4309_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12938$4310_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12941$4311_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12944$4312_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12947$4313_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1295$429_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12950$4314_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12953$4315_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12956$4316_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12959$4317_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12962$4318_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12965$4319_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12968$4320_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12971$4321_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12974$4322_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12977$4323_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1298$430_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12980$4324_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12983$4325_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12986$4326_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12989$4327_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12992$4328_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12995$4329_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:12998$4330_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13001$4331_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13004$4332_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13007$4333_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1301$431_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13010$4334_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13013$4335_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13016$4336_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13019$4337_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13022$4338_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13025$4339_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13028$4340_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13031$4341_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13034$4342_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13037$4343_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1304$432_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13040$4344_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13043$4345_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13046$4346_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13049$4347_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13052$4348_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13055$4349_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13058$4350_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13061$4351_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13064$4352_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13067$4353_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1307$433_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13070$4354_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13073$4355_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13076$4356_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13079$4357_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13082$4358_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13085$4359_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13088$4360_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13091$4361_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13094$4362_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13097$4363_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1310$434_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13100$4364_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13103$4365_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13106$4366_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13109$4367_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13112$4368_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13115$4369_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13118$4370_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13121$4371_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13124$4372_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13127$4373_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1313$435_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13130$4374_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13133$4375_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13136$4376_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13139$4377_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13142$4378_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13145$4379_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13148$4380_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13151$4381_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13154$4382_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13157$4383_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1316$436_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13160$4384_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13163$4385_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13166$4386_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13169$4387_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13172$4388_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13175$4389_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13178$4390_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13181$4391_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13184$4392_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13187$4393_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1319$437_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13190$4394_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13193$4395_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13196$4396_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13199$4397_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13202$4398_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13205$4399_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13208$4400_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13211$4401_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13214$4402_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13217$4403_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1322$438_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13220$4404_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13223$4405_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13226$4406_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13229$4407_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13232$4408_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13235$4409_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13238$4410_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13241$4411_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13244$4412_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13247$4413_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1325$439_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13250$4414_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13253$4415_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13256$4416_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13259$4417_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13262$4418_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13265$4419_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13268$4420_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13271$4421_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13274$4422_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13277$4423_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1328$440_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13280$4424_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13283$4425_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13286$4426_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13289$4427_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13292$4428_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13295$4429_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13298$4430_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13301$4431_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13304$4432_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13307$4433_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1331$441_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13310$4434_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13313$4435_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13316$4436_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13319$4437_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13322$4438_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13325$4439_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13328$4440_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13331$4441_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13334$4442_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13337$4443_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1334$442_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13340$4444_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13343$4445_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13346$4446_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13349$4447_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13352$4448_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13355$4449_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13358$4450_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13361$4451_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13364$4452_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13367$4453_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1337$443_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13370$4454_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13373$4455_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13376$4456_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13379$4457_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13382$4458_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13385$4459_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13388$4460_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13391$4461_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13394$4462_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13397$4463_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1340$444_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13400$4464_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13403$4465_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13406$4466_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13409$4467_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13412$4468_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13415$4469_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13418$4470_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13421$4471_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13424$4472_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13427$4473_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1343$445_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13430$4474_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13433$4475_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13436$4476_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13439$4477_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13442$4478_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13445$4479_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13448$4480_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13451$4481_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13454$4482_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13457$4483_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1346$446_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13460$4484_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13463$4485_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13466$4486_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13469$4487_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13472$4488_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13475$4489_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13478$4490_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13481$4491_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13484$4492_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13487$4493_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1349$447_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13490$4494_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13493$4495_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13496$4496_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13499$4497_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13502$4498_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13505$4499_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13508$4500_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13511$4501_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13514$4502_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13517$4503_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1352$448_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13520$4504_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13523$4505_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13526$4506_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13529$4507_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13532$4508_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13535$4509_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13538$4510_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13541$4511_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13544$4512_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13547$4513_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1355$449_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13550$4514_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13553$4515_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13556$4516_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13559$4517_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13562$4518_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13565$4519_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13568$4520_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13571$4521_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13574$4522_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13577$4523_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1358$450_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13580$4524_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13583$4525_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13586$4526_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13589$4527_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13592$4528_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13595$4529_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13598$4530_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13601$4531_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13604$4532_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13607$4533_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1361$451_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13610$4534_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13613$4535_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13616$4536_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13619$4537_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13622$4538_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13625$4539_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13628$4540_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13631$4541_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13634$4542_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13637$4543_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1364$452_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13640$4544_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13643$4545_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13646$4546_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13649$4547_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13652$4548_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13655$4549_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13658$4550_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13661$4551_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13664$4552_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13667$4553_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1367$453_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13670$4554_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13673$4555_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13676$4556_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13679$4557_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13682$4558_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13685$4559_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13688$4560_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13691$4561_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13694$4562_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13697$4563_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1370$454_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13700$4564_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13703$4565_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13706$4566_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13709$4567_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13712$4568_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13715$4569_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13718$4570_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13721$4571_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13724$4572_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13727$4573_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1373$455_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13730$4574_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13733$4575_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13736$4576_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13739$4577_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13742$4578_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13745$4579_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13748$4580_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13751$4581_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13754$4582_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13757$4583_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1376$456_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13760$4584_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13763$4585_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13766$4586_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13769$4587_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13772$4588_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13775$4589_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13778$4590_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13781$4591_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13784$4592_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13787$4593_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1379$457_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13790$4594_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13793$4595_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13796$4596_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13799$4597_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13802$4598_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13805$4599_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13808$4600_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13811$4601_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13814$4602_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13817$4603_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1382$458_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13820$4604_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13823$4605_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13826$4606_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13829$4607_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13832$4608_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13835$4609_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13838$4610_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13841$4611_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13844$4612_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13847$4613_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1385$459_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13850$4614_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13853$4615_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13856$4616_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13859$4617_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13862$4618_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13865$4619_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13868$4620_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13871$4621_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13874$4622_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13877$4623_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1388$460_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13880$4624_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13883$4625_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13886$4626_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13889$4627_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13892$4628_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13895$4629_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13898$4630_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13901$4631_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13904$4632_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13907$4633_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1391$461_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13910$4634_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13913$4635_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13916$4636_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13919$4637_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13922$4638_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13925$4639_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13928$4640_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13931$4641_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13934$4642_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13937$4643_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1394$462_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13940$4644_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13943$4645_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13946$4646_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13949$4647_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13952$4648_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13955$4649_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13958$4650_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13961$4651_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13964$4652_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13967$4653_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1397$463_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13970$4654_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13973$4655_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13976$4656_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13979$4657_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13982$4658_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13985$4659_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13988$4660_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13991$4661_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13994$4662_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:13997$4663_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1400$464_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14000$4664_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14003$4665_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14006$4666_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14009$4667_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14012$4668_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14015$4669_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14018$4670_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14021$4671_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14024$4672_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14027$4673_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1403$465_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14030$4674_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14033$4675_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14036$4676_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14039$4677_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14042$4678_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14045$4679_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14048$4680_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14051$4681_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14054$4682_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14057$4683_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1406$466_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14060$4684_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14063$4685_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14066$4686_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14069$4687_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14072$4688_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14075$4689_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14078$4690_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14081$4691_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14084$4692_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14087$4693_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1409$467_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14090$4694_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14093$4695_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14096$4696_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14099$4697_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14102$4698_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14105$4699_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14108$4700_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14111$4701_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14114$4702_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14117$4703_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1412$468_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14120$4704_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14123$4705_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14126$4706_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14129$4707_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14132$4708_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14135$4709_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14138$4710_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14141$4711_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14144$4712_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14147$4713_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1415$469_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14150$4714_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14153$4715_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14156$4716_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14159$4717_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14162$4718_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14165$4719_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14168$4720_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14171$4721_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14174$4722_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14177$4723_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1418$470_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14180$4724_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14183$4725_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14186$4726_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14189$4727_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14192$4728_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14195$4729_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14198$4730_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14201$4731_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14204$4732_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14207$4733_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1421$471_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14210$4734_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14213$4735_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14216$4736_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14219$4737_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14222$4738_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14225$4739_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14228$4740_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14231$4741_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14234$4742_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14237$4743_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1424$472_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14240$4744_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14243$4745_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14246$4746_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14249$4747_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14252$4748_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14255$4749_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14258$4750_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14261$4751_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14264$4752_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14267$4753_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1427$473_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14270$4754_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14273$4755_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14276$4756_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14279$4757_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14282$4758_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14285$4759_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14288$4760_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14291$4761_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14294$4762_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14297$4763_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1430$474_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14300$4764_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14303$4765_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14306$4766_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14309$4767_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14312$4768_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14315$4769_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14318$4770_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14321$4771_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14324$4772_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14327$4773_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1433$475_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14330$4774_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14333$4775_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14336$4776_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14339$4777_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14342$4778_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14345$4779_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14348$4780_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14351$4781_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14354$4782_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14357$4783_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1436$476_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14360$4784_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14363$4785_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14366$4786_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14369$4787_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14372$4788_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14375$4789_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14378$4790_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14381$4791_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14384$4792_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14387$4793_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1439$477_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14390$4794_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14393$4795_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14396$4796_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14399$4797_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14402$4798_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14405$4799_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14408$4800_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14411$4801_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14414$4802_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14417$4803_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1442$478_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14420$4804_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14423$4805_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14426$4806_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14429$4807_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14432$4808_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14435$4809_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14438$4810_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14441$4811_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14444$4812_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14447$4813_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1445$479_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14450$4814_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14453$4815_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14456$4816_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14459$4817_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14462$4818_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14465$4819_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14468$4820_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14471$4821_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14474$4822_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14477$4823_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1448$480_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14480$4824_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14483$4825_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14486$4826_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14489$4827_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14492$4828_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14495$4829_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14498$4830_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14501$4831_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14504$4832_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14507$4833_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1451$481_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14510$4834_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14513$4835_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14516$4836_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14519$4837_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14522$4838_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14525$4839_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14528$4840_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14531$4841_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14534$4842_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14537$4843_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1454$482_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14540$4844_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14543$4845_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14546$4846_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14549$4847_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14552$4848_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14555$4849_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14558$4850_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14561$4851_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14564$4852_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14567$4853_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1457$483_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14570$4854_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14573$4855_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14576$4856_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14579$4857_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14582$4858_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14585$4859_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14588$4860_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14591$4861_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14594$4862_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14597$4863_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1460$484_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14600$4864_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14603$4865_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14606$4866_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14609$4867_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14612$4868_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14615$4869_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14618$4870_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14621$4871_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14624$4872_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14627$4873_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1463$485_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14630$4874_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14633$4875_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14636$4876_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14639$4877_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14642$4878_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14645$4879_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14648$4880_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14651$4881_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14654$4882_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14657$4883_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1466$486_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14660$4884_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14663$4885_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14666$4886_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14669$4887_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14672$4888_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14675$4889_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14678$4890_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14681$4891_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14684$4892_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14687$4893_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1469$487_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14690$4894_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14693$4895_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14696$4896_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14699$4897_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14702$4898_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14705$4899_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14708$4900_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14711$4901_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14714$4902_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14717$4903_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1472$488_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14720$4904_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14723$4905_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14726$4906_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14729$4907_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14732$4908_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14735$4909_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14738$4910_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14741$4911_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14744$4912_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14747$4913_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1475$489_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14750$4914_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14753$4915_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14756$4916_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14759$4917_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14762$4918_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14765$4919_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14768$4920_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14771$4921_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14774$4922_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14777$4923_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1478$490_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14780$4924_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14783$4925_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14786$4926_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14789$4927_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14792$4928_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14795$4929_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14798$4930_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14801$4931_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14804$4932_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14807$4933_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1481$491_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14810$4934_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14813$4935_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14816$4936_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14819$4937_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14822$4938_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14825$4939_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14828$4940_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14831$4941_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14834$4942_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14837$4943_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1484$492_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14840$4944_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14843$4945_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14846$4946_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14849$4947_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14852$4948_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14855$4949_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14858$4950_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14861$4951_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14864$4952_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14867$4953_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1487$493_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14870$4954_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14873$4955_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14876$4956_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14879$4957_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14882$4958_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14885$4959_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14888$4960_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14891$4961_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14894$4962_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14897$4963_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1490$494_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14900$4964_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14903$4965_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14906$4966_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14909$4967_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14912$4968_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14915$4969_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14918$4970_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14921$4971_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14924$4972_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14927$4973_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1493$495_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14930$4974_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14933$4975_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14936$4976_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14939$4977_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14942$4978_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14945$4979_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14948$4980_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14951$4981_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14954$4982_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14957$4983_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1496$496_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14960$4984_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14963$4985_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14966$4986_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14969$4987_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14972$4988_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14975$4989_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14978$4990_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14981$4991_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14984$4992_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14987$4993_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1499$497_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14990$4994_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14993$4995_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14996$4996_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:14999$4997_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15002$4998_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15005$4999_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15008$5000_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15011$5001_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15014$5002_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15017$5003_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1502$498_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15020$5004_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15023$5005_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15026$5006_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15029$5007_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15032$5008_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15035$5009_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15038$5010_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15041$5011_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15044$5012_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15047$5013_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1505$499_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15050$5014_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15053$5015_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15056$5016_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15059$5017_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15062$5018_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15065$5019_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15068$5020_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15071$5021_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15074$5022_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15077$5023_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1508$500_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15080$5024_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15083$5025_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15086$5026_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15089$5027_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15092$5028_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15095$5029_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15098$5030_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15101$5031_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15104$5032_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15107$5033_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1511$501_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15110$5034_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15113$5035_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15116$5036_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15119$5037_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15122$5038_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15125$5039_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15128$5040_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15131$5041_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15134$5042_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15137$5043_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1514$502_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15140$5044_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15143$5045_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15146$5046_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15149$5047_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15152$5048_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15155$5049_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15158$5050_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15161$5051_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15164$5052_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15167$5053_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1517$503_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15170$5054_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15173$5055_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15176$5056_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15179$5057_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15182$5058_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15185$5059_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15188$5060_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15191$5061_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15194$5062_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15197$5063_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1520$504_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15200$5064_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15203$5065_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15206$5066_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15209$5067_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15212$5068_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15215$5069_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15218$5070_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15221$5071_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15224$5072_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15227$5073_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1523$505_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15230$5074_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15233$5075_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15236$5076_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15239$5077_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15242$5078_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15245$5079_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15248$5080_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15251$5081_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15254$5082_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15257$5083_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1526$506_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15260$5084_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15263$5085_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15266$5086_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15269$5087_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15272$5088_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15275$5089_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15278$5090_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15281$5091_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15284$5092_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15287$5093_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1529$507_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15290$5094_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15293$5095_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15296$5096_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15299$5097_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15302$5098_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15305$5099_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15308$5100_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15311$5101_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15314$5102_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15317$5103_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1532$508_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15320$5104_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15323$5105_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15326$5106_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15329$5107_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15332$5108_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15335$5109_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15338$5110_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15341$5111_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15344$5112_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15347$5113_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1535$509_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15350$5114_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15353$5115_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15356$5116_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15359$5117_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15362$5118_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15365$5119_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15368$5120_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15371$5121_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15374$5122_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15377$5123_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1538$510_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15380$5124_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15383$5125_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15386$5126_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15389$5127_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15392$5128_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15395$5129_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15398$5130_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15401$5131_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15404$5132_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15407$5133_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1541$511_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15410$5134_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15413$5135_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15416$5136_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15419$5137_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15422$5138_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15425$5139_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15428$5140_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15431$5141_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15434$5142_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15437$5143_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1544$512_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15440$5144_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15443$5145_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15446$5146_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15449$5147_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15452$5148_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15455$5149_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15458$5150_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15461$5151_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15464$5152_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15467$5153_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1547$513_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15470$5154_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15473$5155_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15476$5156_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15479$5157_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15482$5158_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15485$5159_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15488$5160_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15491$5161_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15494$5162_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15497$5163_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1550$514_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15500$5164_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15503$5165_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15506$5166_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15509$5167_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15512$5168_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15515$5169_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15518$5170_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15521$5171_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15524$5172_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15527$5173_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1553$515_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15530$5174_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15533$5175_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15536$5176_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15539$5177_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15542$5178_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15545$5179_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15548$5180_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15551$5181_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15554$5182_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15557$5183_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1556$516_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15560$5184_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15563$5185_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15566$5186_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15569$5187_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15572$5188_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15575$5189_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15578$5190_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15581$5191_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15584$5192_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15587$5193_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1559$517_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15590$5194_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15593$5195_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15596$5196_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15599$5197_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15602$5198_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15605$5199_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15608$5200_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15611$5201_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15614$5202_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15617$5203_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1562$518_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15620$5204_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15623$5205_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15626$5206_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15629$5207_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15632$5208_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15635$5209_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15638$5210_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15641$5211_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15644$5212_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15647$5213_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1565$519_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15650$5214_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15653$5215_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15656$5216_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15659$5217_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15662$5218_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15665$5219_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15668$5220_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15671$5221_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15674$5222_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15677$5223_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1568$520_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15680$5224_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15683$5225_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15686$5226_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15689$5227_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15692$5228_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15695$5229_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15698$5230_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15701$5231_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15704$5232_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15707$5233_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1571$521_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15710$5234_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15713$5235_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15716$5236_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15719$5237_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15722$5238_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15725$5239_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15728$5240_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15731$5241_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15734$5242_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15737$5243_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1574$522_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15740$5244_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15743$5245_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15746$5246_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15749$5247_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15752$5248_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15755$5249_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15758$5250_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15761$5251_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15764$5252_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15767$5253_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1577$523_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15770$5254_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15773$5255_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15776$5256_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15779$5257_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15782$5258_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15785$5259_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15788$5260_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15791$5261_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15794$5262_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15797$5263_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1580$524_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15800$5264_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15803$5265_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15806$5266_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15809$5267_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15812$5268_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15815$5269_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15818$5270_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15821$5271_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15824$5272_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15827$5273_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1583$525_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15830$5274_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15833$5275_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15836$5276_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15839$5277_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15842$5278_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15845$5279_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15848$5280_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15851$5281_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15854$5282_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15857$5283_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1586$526_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15860$5284_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15863$5285_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15866$5286_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15869$5287_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15872$5288_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15875$5289_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15878$5290_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15881$5291_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15884$5292_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15887$5293_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1589$527_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15890$5294_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15893$5295_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15896$5296_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15899$5297_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15902$5298_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15905$5299_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15908$5300_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15911$5301_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15914$5302_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15917$5303_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1592$528_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15920$5304_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15923$5305_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15926$5306_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15929$5307_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15932$5308_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15935$5309_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15938$5310_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15941$5311_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15944$5312_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15947$5313_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1595$529_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15950$5314_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15953$5315_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15956$5316_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15959$5317_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15962$5318_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15965$5319_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15968$5320_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15971$5321_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15974$5322_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15977$5323_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1598$530_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15980$5324_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15983$5325_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15986$5326_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15989$5327_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15992$5328_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15995$5329_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:15998$5330_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16001$5331_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16004$5332_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16007$5333_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1601$531_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16010$5334_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16013$5335_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16016$5336_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16019$5337_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16022$5338_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16025$5339_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16028$5340_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16031$5341_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16034$5342_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16037$5343_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1604$532_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16040$5344_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16043$5345_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16046$5346_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16049$5347_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16052$5348_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16055$5349_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16058$5350_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16061$5351_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16064$5352_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16067$5353_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1607$533_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16070$5354_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16073$5355_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16076$5356_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16079$5357_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16082$5358_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16085$5359_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16088$5360_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16091$5361_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16094$5362_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16097$5363_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1610$534_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16100$5364_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16103$5365_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16106$5366_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16109$5367_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16112$5368_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16115$5369_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16118$5370_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16121$5371_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16124$5372_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16127$5373_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1613$535_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16130$5374_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16133$5375_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16136$5376_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16139$5377_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16142$5378_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16145$5379_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16148$5380_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16151$5381_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16154$5382_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16157$5383_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1616$536_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16160$5384_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16163$5385_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16166$5386_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16169$5387_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16172$5388_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16175$5389_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16178$5390_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16181$5391_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16184$5392_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16187$5393_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1619$537_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16190$5394_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16193$5395_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16196$5396_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16199$5397_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16202$5398_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16205$5399_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16208$5400_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16211$5401_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16214$5402_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16217$5403_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1622$538_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16220$5404_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16223$5405_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16226$5406_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16229$5407_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16232$5408_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16235$5409_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16238$5410_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16241$5411_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16244$5412_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16247$5413_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1625$539_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16250$5414_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16253$5415_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16256$5416_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16259$5417_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16262$5418_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16265$5419_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16268$5420_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16271$5421_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16274$5422_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16277$5423_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1628$540_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16280$5424_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16283$5425_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16286$5426_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16289$5427_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16292$5428_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16295$5429_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16298$5430_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16301$5431_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16304$5432_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16307$5433_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1631$541_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16310$5434_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16313$5435_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16316$5436_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16319$5437_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16322$5438_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16325$5439_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16328$5440_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16331$5441_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16334$5442_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16337$5443_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1634$542_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16340$5444_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16343$5445_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16346$5446_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16349$5447_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16352$5448_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16355$5449_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16358$5450_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16361$5451_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16364$5452_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16367$5453_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1637$543_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16370$5454_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16373$5455_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16376$5456_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16379$5457_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16382$5458_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16385$5459_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16388$5460_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16391$5461_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16394$5462_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16397$5463_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1640$544_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16400$5464_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16403$5465_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16406$5466_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16409$5467_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16412$5468_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16415$5469_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16418$5470_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16421$5471_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16424$5472_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16427$5473_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1643$545_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16430$5474_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16433$5475_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16436$5476_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16439$5477_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16442$5478_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16445$5479_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16448$5480_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16451$5481_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16454$5482_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16457$5483_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1646$546_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16460$5484_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16463$5485_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16466$5486_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16469$5487_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16472$5488_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16475$5489_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16478$5490_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16481$5491_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16484$5492_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16487$5493_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1649$547_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16490$5494_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16493$5495_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16496$5496_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16499$5497_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16502$5498_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16505$5499_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16508$5500_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16511$5501_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16514$5502_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16517$5503_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1652$548_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16520$5504_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16523$5505_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16526$5506_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16529$5507_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16532$5508_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16535$5509_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16538$5510_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16541$5511_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16544$5512_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16547$5513_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1655$549_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16550$5514_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16553$5515_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16556$5516_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16559$5517_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16562$5518_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16565$5519_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16568$5520_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16571$5521_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16574$5522_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16577$5523_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1658$550_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16580$5524_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16583$5525_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16586$5526_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16589$5527_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16592$5528_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16595$5529_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16598$5530_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16601$5531_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16604$5532_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16607$5533_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1661$551_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16610$5534_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16613$5535_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16616$5536_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16619$5537_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16622$5538_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16625$5539_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16628$5540_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16631$5541_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16634$5542_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16637$5543_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1664$552_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16640$5544_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16643$5545_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16646$5546_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16649$5547_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16652$5548_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16655$5549_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16658$5550_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16661$5551_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16664$5552_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16667$5553_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1667$553_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16670$5554_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16673$5555_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16676$5556_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16679$5557_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16682$5558_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16685$5559_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16688$5560_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16691$5561_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16694$5562_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16697$5563_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1670$554_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16700$5564_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16703$5565_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16706$5566_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16709$5567_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16712$5568_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16715$5569_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16718$5570_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16721$5571_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16724$5572_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16727$5573_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1673$555_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16730$5574_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16733$5575_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16736$5576_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16739$5577_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16742$5578_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16745$5579_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16748$5580_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16751$5581_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16754$5582_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16757$5583_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1676$556_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16760$5584_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16763$5585_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16766$5586_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16769$5587_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16772$5588_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16775$5589_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16778$5590_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16781$5591_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16784$5592_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16787$5593_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1679$557_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16790$5594_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16793$5595_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16796$5596_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16799$5597_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16802$5598_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16805$5599_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16808$5600_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16811$5601_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16814$5602_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16817$5603_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1682$558_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16820$5604_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16823$5605_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16826$5606_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16829$5607_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16832$5608_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16835$5609_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16838$5610_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16841$5611_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16844$5612_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16847$5613_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1685$559_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16850$5614_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16853$5615_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16856$5616_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16859$5617_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16862$5618_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16865$5619_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16868$5620_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16871$5621_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16874$5622_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16877$5623_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1688$560_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16880$5624_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16883$5625_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16886$5626_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16889$5627_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16892$5628_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16895$5629_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16898$5630_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16901$5631_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16904$5632_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16907$5633_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1691$561_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16910$5634_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16913$5635_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16916$5636_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16919$5637_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16922$5638_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16925$5639_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16928$5640_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16931$5641_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16934$5642_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16937$5643_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1694$562_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16940$5644_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16943$5645_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16946$5646_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16949$5647_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16952$5648_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16955$5649_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16958$5650_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16961$5651_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16964$5652_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16967$5653_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1697$563_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16970$5654_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16973$5655_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16976$5656_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16979$5657_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16982$5658_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16985$5659_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16988$5660_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16991$5661_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16994$5662_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:16997$5663_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1700$564_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17000$5664_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17003$5665_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17006$5666_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17009$5667_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17012$5668_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17015$5669_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17018$5670_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17021$5671_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17024$5672_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17027$5673_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1703$565_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17030$5674_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17033$5675_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17036$5676_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17039$5677_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17042$5678_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17045$5679_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17048$5680_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17051$5681_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17054$5682_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17057$5683_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1706$566_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17060$5684_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17063$5685_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17066$5686_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17069$5687_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17072$5688_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17075$5689_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17078$5690_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17081$5691_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17084$5692_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17087$5693_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1709$567_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17090$5694_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17093$5695_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17096$5696_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17099$5697_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17102$5698_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17105$5699_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17108$5700_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17111$5701_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17114$5702_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17117$5703_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1712$568_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17120$5704_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17123$5705_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17126$5706_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17129$5707_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17132$5708_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17135$5709_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17138$5710_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17141$5711_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17144$5712_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17147$5713_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1715$569_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17150$5714_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17153$5715_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17156$5716_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17159$5717_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17162$5718_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17165$5719_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17168$5720_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17171$5721_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17174$5722_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17177$5723_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1718$570_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17180$5724_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17183$5725_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17186$5726_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17189$5727_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17192$5728_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17195$5729_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17198$5730_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17201$5731_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17204$5732_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17207$5733_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1721$571_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17210$5734_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17213$5735_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17216$5736_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17219$5737_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17222$5738_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17225$5739_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17228$5740_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17231$5741_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17234$5742_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17237$5743_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1724$572_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17240$5744_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17243$5745_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17246$5746_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17249$5747_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17252$5748_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17255$5749_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17258$5750_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17261$5751_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17264$5752_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17267$5753_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1727$573_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17270$5754_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17273$5755_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17276$5756_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17279$5757_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17282$5758_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17285$5759_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17288$5760_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17291$5761_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17294$5762_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17297$5763_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1730$574_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17300$5764_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17303$5765_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17306$5766_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17309$5767_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17312$5768_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17315$5769_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17318$5770_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17321$5771_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17324$5772_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17327$5773_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1733$575_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17330$5774_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17333$5775_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17336$5776_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17339$5777_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17342$5778_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17345$5779_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17348$5780_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17351$5781_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17354$5782_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17357$5783_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1736$576_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17360$5784_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17363$5785_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17366$5786_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17369$5787_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17372$5788_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17375$5789_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17378$5790_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17381$5791_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17384$5792_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17387$5793_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1739$577_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17390$5794_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17393$5795_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17396$5796_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17399$5797_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17402$5798_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17405$5799_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17408$5800_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17411$5801_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17414$5802_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17417$5803_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1742$578_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17420$5804_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17423$5805_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17426$5806_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17429$5807_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17432$5808_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17435$5809_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17438$5810_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17441$5811_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17444$5812_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17447$5813_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1745$579_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17450$5814_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17453$5815_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17456$5816_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17459$5817_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17462$5818_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17465$5819_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17468$5820_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17471$5821_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17474$5822_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17477$5823_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1748$580_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17480$5824_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17483$5825_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17486$5826_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17489$5827_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17492$5828_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17495$5829_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17498$5830_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17501$5831_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17504$5832_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17507$5833_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1751$581_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17510$5834_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17513$5835_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17516$5836_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17519$5837_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17522$5838_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17525$5839_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17528$5840_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17531$5841_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17534$5842_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17537$5843_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1754$582_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17540$5844_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17543$5845_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17546$5846_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17549$5847_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17552$5848_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17555$5849_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17558$5850_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17561$5851_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17564$5852_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17567$5853_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1757$583_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17570$5854_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17573$5855_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17576$5856_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17579$5857_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17582$5858_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17585$5859_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17588$5860_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17591$5861_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17594$5862_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17597$5863_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1760$584_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17600$5864_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17603$5865_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17606$5866_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17609$5867_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17612$5868_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17615$5869_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17618$5870_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17621$5871_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17624$5872_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17627$5873_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1763$585_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17630$5874_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17633$5875_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17636$5876_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17639$5877_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17642$5878_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17645$5879_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17648$5880_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17651$5881_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17654$5882_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17657$5883_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1766$586_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17660$5884_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17663$5885_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17666$5886_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17669$5887_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17672$5888_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17675$5889_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17678$5890_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17681$5891_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17684$5892_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17687$5893_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1769$587_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17690$5894_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17693$5895_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17696$5896_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17699$5897_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17702$5898_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17705$5899_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17708$5900_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17711$5901_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17714$5902_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17717$5903_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1772$588_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17720$5904_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17723$5905_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17726$5906_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17729$5907_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17732$5908_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17735$5909_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17738$5910_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17741$5911_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17744$5912_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17747$5913_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1775$589_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17750$5914_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17753$5915_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17756$5916_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17759$5917_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17762$5918_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17765$5919_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17768$5920_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17771$5921_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17774$5922_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17777$5923_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1778$590_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17780$5924_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17783$5925_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17786$5926_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17789$5927_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17792$5928_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17795$5929_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17798$5930_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17801$5931_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17804$5932_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17807$5933_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1781$591_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17810$5934_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17813$5935_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17816$5936_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17819$5937_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17822$5938_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17825$5939_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17828$5940_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17831$5941_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17834$5942_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17837$5943_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1784$592_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17840$5944_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17843$5945_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17846$5946_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17849$5947_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17852$5948_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17855$5949_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17858$5950_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17861$5951_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17864$5952_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17867$5953_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1787$593_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17870$5954_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17873$5955_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17876$5956_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17879$5957_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17882$5958_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17885$5959_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17888$5960_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17891$5961_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17894$5962_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17897$5963_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1790$594_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17900$5964_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17903$5965_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17906$5966_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17909$5967_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17912$5968_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17915$5969_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17918$5970_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17921$5971_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17924$5972_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17927$5973_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1793$595_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17930$5974_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17933$5975_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17936$5976_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17939$5977_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17942$5978_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17945$5979_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17948$5980_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17951$5981_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17954$5982_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17957$5983_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1796$596_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17960$5984_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17963$5985_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17966$5986_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17969$5987_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17972$5988_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17975$5989_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17978$5990_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17981$5991_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17984$5992_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17987$5993_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1799$597_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17990$5994_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17993$5995_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17996$5996_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:17999$5997_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18002$5998_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18005$5999_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18008$6000_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18011$6001_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18014$6002_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18017$6003_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1802$598_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18020$6004_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18023$6005_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18026$6006_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18029$6007_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18032$6008_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18035$6009_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18038$6010_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18041$6011_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18044$6012_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18047$6013_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1805$599_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18050$6014_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18053$6015_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18056$6016_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18059$6017_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18062$6018_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18065$6019_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18068$6020_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18071$6021_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18074$6022_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18077$6023_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1808$600_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18080$6024_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18083$6025_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18086$6026_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18089$6027_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18092$6028_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18095$6029_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18098$6030_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18101$6031_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18104$6032_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18107$6033_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1811$601_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18110$6034_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18113$6035_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18116$6036_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18119$6037_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18122$6038_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18125$6039_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18128$6040_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18131$6041_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18134$6042_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18137$6043_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1814$602_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18140$6044_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18143$6045_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18146$6046_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18149$6047_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18152$6048_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18155$6049_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18158$6050_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18161$6051_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18164$6052_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18167$6053_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1817$603_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18170$6054_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18173$6055_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18176$6056_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18179$6057_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18182$6058_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18185$6059_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18188$6060_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18191$6061_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18194$6062_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18197$6063_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1820$604_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18200$6064_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18203$6065_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18206$6066_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18209$6067_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18212$6068_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18215$6069_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18218$6070_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18221$6071_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18224$6072_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18227$6073_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1823$605_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18230$6074_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18233$6075_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18236$6076_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18239$6077_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18242$6078_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18245$6079_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18248$6080_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18251$6081_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18254$6082_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18257$6083_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1826$606_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18260$6084_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18263$6085_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18266$6086_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18269$6087_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18272$6088_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18275$6089_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18278$6090_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18281$6091_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18284$6092_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18287$6093_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1829$607_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18290$6094_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18293$6095_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18296$6096_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18299$6097_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18302$6098_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18305$6099_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18308$6100_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18311$6101_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18314$6102_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18317$6103_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1832$608_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18320$6104_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18323$6105_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18326$6106_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18329$6107_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18332$6108_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18335$6109_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18338$6110_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18341$6111_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18344$6112_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18347$6113_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1835$609_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18350$6114_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18353$6115_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18356$6116_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18359$6117_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18362$6118_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18365$6119_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18368$6120_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18371$6121_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18374$6122_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18377$6123_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1838$610_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18380$6124_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18383$6125_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18386$6126_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18389$6127_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18392$6128_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18395$6129_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18398$6130_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18401$6131_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18404$6132_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18407$6133_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1841$611_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18410$6134_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18413$6135_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18416$6136_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18419$6137_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18422$6138_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18425$6139_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18428$6140_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18431$6141_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18434$6142_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18437$6143_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1844$612_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18440$6144_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18443$6145_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18446$6146_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18449$6147_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18452$6148_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18455$6149_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18458$6150_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18461$6151_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18464$6152_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18467$6153_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1847$613_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18470$6154_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18473$6155_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18476$6156_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18479$6157_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18482$6158_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18485$6159_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18488$6160_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18491$6161_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18494$6162_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18497$6163_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1850$614_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18500$6164_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18503$6165_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18506$6166_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18509$6167_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18512$6168_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18515$6169_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18518$6170_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18521$6171_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18524$6172_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18527$6173_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1853$615_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18530$6174_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18533$6175_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18536$6176_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18539$6177_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18542$6178_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18545$6179_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18548$6180_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18551$6181_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18554$6182_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18557$6183_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1856$616_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18560$6184_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18563$6185_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18566$6186_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18569$6187_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18572$6188_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18575$6189_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18578$6190_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18581$6191_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18584$6192_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18587$6193_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1859$617_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18590$6194_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18593$6195_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18596$6196_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18599$6197_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18602$6198_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18605$6199_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18608$6200_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18611$6201_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18614$6202_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18617$6203_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1862$618_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18620$6204_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18623$6205_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18626$6206_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18629$6207_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18632$6208_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18635$6209_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18638$6210_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18641$6211_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18644$6212_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18647$6213_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1865$619_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18650$6214_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18653$6215_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18656$6216_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18659$6217_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18662$6218_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18665$6219_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18668$6220_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18671$6221_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18674$6222_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18677$6223_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1868$620_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18680$6224_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18683$6225_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18686$6226_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18689$6227_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18692$6228_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18695$6229_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18698$6230_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18701$6231_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18704$6232_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18707$6233_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1871$621_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18710$6234_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18713$6235_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18716$6236_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18719$6237_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18722$6238_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18725$6239_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18728$6240_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18731$6241_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18734$6242_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18737$6243_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1874$622_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18740$6244_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18743$6245_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18746$6246_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18749$6247_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18752$6248_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18755$6249_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18758$6250_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18761$6251_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18764$6252_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18767$6253_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1877$623_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18770$6254_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18773$6255_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18776$6256_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18779$6257_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18782$6258_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18785$6259_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18788$6260_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18791$6261_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18794$6262_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18797$6263_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1880$624_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18800$6264_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18803$6265_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18806$6266_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18809$6267_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18812$6268_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18815$6269_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18818$6270_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18821$6271_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18824$6272_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18827$6273_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1883$625_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18830$6274_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18833$6275_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18836$6276_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18839$6277_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18842$6278_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18845$6279_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18848$6280_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18851$6281_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18854$6282_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18857$6283_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1886$626_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18860$6284_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18863$6285_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18866$6286_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18869$6287_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18872$6288_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18875$6289_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18878$6290_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18881$6291_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18884$6292_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18887$6293_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1889$627_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18890$6294_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18893$6295_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18896$6296_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18899$6297_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18902$6298_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:18905$6299_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1892$628_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1895$629_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1898$630_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1901$631_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1904$632_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1907$633_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1910$634_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1913$635_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1916$636_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1919$637_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1922$638_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1925$639_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1928$640_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1931$641_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1934$642_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1937$643_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1940$644_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1943$645_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1946$646_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1949$647_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1952$648_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1955$649_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1958$650_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1961$651_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1964$652_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1967$653_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1970$654_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1973$655_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1976$656_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1979$657_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1982$658_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1985$659_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1988$660_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1991$661_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1994$662_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:1997$663_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2000$664_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2003$665_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2006$666_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2009$667_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2012$668_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2015$669_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2018$670_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2021$671_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2024$672_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2027$673_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2030$674_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2033$675_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2036$676_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2039$677_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2042$678_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2045$679_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2048$680_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2051$681_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2054$682_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2057$683_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2060$684_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2063$685_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2066$686_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2069$687_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2072$688_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2075$689_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2078$690_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2081$691_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2084$692_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2087$693_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2090$694_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2093$695_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2096$696_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2099$697_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2102$698_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2105$699_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2108$700_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2111$701_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2114$702_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2117$703_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2120$704_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2123$705_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2126$706_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2129$707_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2132$708_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2135$709_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2138$710_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2141$711_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2144$712_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2147$713_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2150$714_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2153$715_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2156$716_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2159$717_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2162$718_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2165$719_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2168$720_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2171$721_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2174$722_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2177$723_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2180$724_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2183$725_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2186$726_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2189$727_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2192$728_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2195$729_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2198$730_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2201$731_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2204$732_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2207$733_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2210$734_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2213$735_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2216$736_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2219$737_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2222$738_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2225$739_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2228$740_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2231$741_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2234$742_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2237$743_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2240$744_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2243$745_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2246$746_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2249$747_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2252$748_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2255$749_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2258$750_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2261$751_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2264$752_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2267$753_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2270$754_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2273$755_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2276$756_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2279$757_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2282$758_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2285$759_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2288$760_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2291$761_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2294$762_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2297$763_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2300$764_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2303$765_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2306$766_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2309$767_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2312$768_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2315$769_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2318$770_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2321$771_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2324$772_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2327$773_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2330$774_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2333$775_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2336$776_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2339$777_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2342$778_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2345$779_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2348$780_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2351$781_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2354$782_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2357$783_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2360$784_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2363$785_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2366$786_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2369$787_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2372$788_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2375$789_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2378$790_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2381$791_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2384$792_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2387$793_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2390$794_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2393$795_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2396$796_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2399$797_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2402$798_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2405$799_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2408$800_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2411$801_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2414$802_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2417$803_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2420$804_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2423$805_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2426$806_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2429$807_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2432$808_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2435$809_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2438$810_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2441$811_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2444$812_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2447$813_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2450$814_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2453$815_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2456$816_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2459$817_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2462$818_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2465$819_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2468$820_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2471$821_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2474$822_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2477$823_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2480$824_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2483$825_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2486$826_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2489$827_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2492$828_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2495$829_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2498$830_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2501$831_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2504$832_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2507$833_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2510$834_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2513$835_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2516$836_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2519$837_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2522$838_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2525$839_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2528$840_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2531$841_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2534$842_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2537$843_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2540$844_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2543$845_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2546$846_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2549$847_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2552$848_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2555$849_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2558$850_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2561$851_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2564$852_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2567$853_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2570$854_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2573$855_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2576$856_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2579$857_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2582$858_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2585$859_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2588$860_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2591$861_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2594$862_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2597$863_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2600$864_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2603$865_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2606$866_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2609$867_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2612$868_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2615$869_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2618$870_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2621$871_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2624$872_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2627$873_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2630$874_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2633$875_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2636$876_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2639$877_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2642$878_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2645$879_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2648$880_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2651$881_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2654$882_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2657$883_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2660$884_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2663$885_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2666$886_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2669$887_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2672$888_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2675$889_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2678$890_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2681$891_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2684$892_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2687$893_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2690$894_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2693$895_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2696$896_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2699$897_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2702$898_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2705$899_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2708$900_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2711$901_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2714$902_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2717$903_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2720$904_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2723$905_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2726$906_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2729$907_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2732$908_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2735$909_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2738$910_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2741$911_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2744$912_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2747$913_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2750$914_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2753$915_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2756$916_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2759$917_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2762$918_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2765$919_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2768$920_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2771$921_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2774$922_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2777$923_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2780$924_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2783$925_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2786$926_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2789$927_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2792$928_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2795$929_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2798$930_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2801$931_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2804$932_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2807$933_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2810$934_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2813$935_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2816$936_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2819$937_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2822$938_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2825$939_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2828$940_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2831$941_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2834$942_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2837$943_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2840$944_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2843$945_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2846$946_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2849$947_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2852$948_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2855$949_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2858$950_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2861$951_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2864$952_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2867$953_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2870$954_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2873$955_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2876$956_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2879$957_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2882$958_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2885$959_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2888$960_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2891$961_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2894$962_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2897$963_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2900$964_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2903$965_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2906$966_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2909$967_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2912$968_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2915$969_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2918$970_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2921$971_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2924$972_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2927$973_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2930$974_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2933$975_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2936$976_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2939$977_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2942$978_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2945$979_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2948$980_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2951$981_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2954$982_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2957$983_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2960$984_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2963$985_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2966$986_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2969$987_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2972$988_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2975$989_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2978$990_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2981$991_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2984$992_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2987$993_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2990$994_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2993$995_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2996$996_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:2999$997_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3002$998_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3005$999_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3008$1000_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3011$1001_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3014$1002_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3017$1003_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3020$1004_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3023$1005_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3026$1006_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3029$1007_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3032$1008_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3035$1009_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3038$1010_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3041$1011_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3044$1012_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3047$1013_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3050$1014_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3053$1015_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3056$1016_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3059$1017_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3062$1018_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3065$1019_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3068$1020_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3071$1021_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3074$1022_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3077$1023_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3080$1024_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3083$1025_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3086$1026_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3089$1027_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3092$1028_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3095$1029_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3098$1030_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3101$1031_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3104$1032_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3107$1033_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3110$1034_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3113$1035_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3116$1036_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3119$1037_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3122$1038_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3125$1039_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3128$1040_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3131$1041_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3134$1042_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3137$1043_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3140$1044_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3143$1045_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3146$1046_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3149$1047_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3152$1048_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3155$1049_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3158$1050_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3161$1051_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3164$1052_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3167$1053_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3170$1054_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3173$1055_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3176$1056_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3179$1057_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3182$1058_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3185$1059_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3188$1060_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3191$1061_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3194$1062_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3197$1063_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:320$104_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:320$104_EN  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3200$1064_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3203$1065_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3206$1066_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3209$1067_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3212$1068_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3215$1069_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3218$1070_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3221$1071_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3224$1072_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3227$1073_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:323$105_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3230$1074_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3233$1075_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3236$1076_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3239$1077_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3242$1078_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3245$1079_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3248$1080_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3251$1081_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3254$1082_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3257$1083_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:326$106_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3260$1084_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3263$1085_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3266$1086_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3269$1087_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3272$1088_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3275$1089_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3278$1090_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3281$1091_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3284$1092_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3287$1093_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:329$107_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3290$1094_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3293$1095_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3296$1096_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3299$1097_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3302$1098_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3305$1099_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3308$1100_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3311$1101_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3314$1102_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3317$1103_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:332$108_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3320$1104_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3323$1105_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3326$1106_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3329$1107_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3332$1108_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3335$1109_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3338$1110_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3341$1111_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3344$1112_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3347$1113_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:335$109_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3350$1114_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3353$1115_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3356$1116_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3359$1117_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3362$1118_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3365$1119_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3368$1120_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3371$1121_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3374$1122_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3377$1123_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:338$110_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3380$1124_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3383$1125_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3386$1126_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3389$1127_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3392$1128_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3395$1129_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3398$1130_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3401$1131_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3404$1132_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3407$1133_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:341$111_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3410$1134_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3413$1135_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3416$1136_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3419$1137_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3422$1138_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3425$1139_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3428$1140_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3431$1141_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3434$1142_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3437$1143_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:344$112_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3440$1144_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3443$1145_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3446$1146_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3449$1147_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3452$1148_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3455$1149_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3458$1150_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3461$1151_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3464$1152_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3467$1153_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:347$113_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3470$1154_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3473$1155_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3476$1156_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3479$1157_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3482$1158_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3485$1159_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3488$1160_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3491$1161_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3494$1162_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3497$1163_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:350$114_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3500$1164_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3503$1165_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3506$1166_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3509$1167_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3512$1168_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3515$1169_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3518$1170_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3521$1171_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3524$1172_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3527$1173_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:353$115_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3530$1174_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3533$1175_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3536$1176_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3539$1177_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3542$1178_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3545$1179_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3548$1180_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3551$1181_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3554$1182_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3557$1183_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:356$116_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3560$1184_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3563$1185_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3566$1186_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3569$1187_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3572$1188_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3575$1189_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3578$1190_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3581$1191_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3584$1192_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3587$1193_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:359$117_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3590$1194_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3593$1195_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3596$1196_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3599$1197_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3602$1198_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3605$1199_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3608$1200_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3611$1201_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3614$1202_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3617$1203_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:362$118_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3620$1204_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3623$1205_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3626$1206_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3629$1207_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3632$1208_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3635$1209_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3638$1210_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3641$1211_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3644$1212_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3647$1213_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:365$119_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3650$1214_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3653$1215_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3656$1216_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3659$1217_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3662$1218_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3665$1219_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3668$1220_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3671$1221_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3674$1222_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3677$1223_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:368$120_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3680$1224_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3683$1225_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3686$1226_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3689$1227_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3692$1228_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3695$1229_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3698$1230_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3701$1231_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3704$1232_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3707$1233_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:371$121_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3710$1234_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3713$1235_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3716$1236_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3719$1237_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3722$1238_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3725$1239_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3728$1240_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3731$1241_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3734$1242_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3737$1243_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:374$122_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3740$1244_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3743$1245_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3746$1246_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3749$1247_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3752$1248_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3755$1249_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3758$1250_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3761$1251_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3764$1252_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3767$1253_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:377$123_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3770$1254_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3773$1255_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3776$1256_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3779$1257_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3782$1258_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3785$1259_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3788$1260_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3791$1261_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3794$1262_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3797$1263_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:380$124_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3800$1264_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3803$1265_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3806$1266_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3809$1267_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3812$1268_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3815$1269_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3818$1270_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3821$1271_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3824$1272_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3827$1273_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:383$125_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3830$1274_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3833$1275_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3836$1276_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3839$1277_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3842$1278_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3845$1279_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3848$1280_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3851$1281_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3854$1282_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3857$1283_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:386$126_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3860$1284_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3863$1285_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3866$1286_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3869$1287_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3872$1288_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3875$1289_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3878$1290_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3881$1291_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3884$1292_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3887$1293_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:389$127_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3890$1294_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3893$1295_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3896$1296_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3899$1297_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3902$1298_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3905$1299_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3908$1300_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3911$1301_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3914$1302_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3917$1303_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:392$128_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3920$1304_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3923$1305_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3926$1306_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3929$1307_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3932$1308_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3935$1309_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3938$1310_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3941$1311_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3944$1312_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3947$1313_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:395$129_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3950$1314_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3953$1315_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3956$1316_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3959$1317_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3962$1318_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3965$1319_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3968$1320_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3971$1321_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3974$1322_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3977$1323_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:398$130_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3980$1324_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3983$1325_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3986$1326_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3989$1327_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3992$1328_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3995$1329_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:3998$1330_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4001$1331_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4004$1332_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4007$1333_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:401$131_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4010$1334_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4013$1335_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4016$1336_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4019$1337_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4022$1338_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4025$1339_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4028$1340_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4031$1341_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4034$1342_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4037$1343_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:404$132_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4040$1344_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4043$1345_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4046$1346_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4049$1347_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4052$1348_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4055$1349_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4058$1350_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4061$1351_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4064$1352_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4067$1353_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:407$133_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4070$1354_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4073$1355_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4076$1356_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4079$1357_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4082$1358_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4085$1359_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4088$1360_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4091$1361_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4094$1362_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4097$1363_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:410$134_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4100$1364_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4103$1365_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4106$1366_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4109$1367_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4112$1368_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4115$1369_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4118$1370_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4121$1371_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4124$1372_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4127$1373_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:413$135_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4130$1374_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4133$1375_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4136$1376_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4139$1377_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4142$1378_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4145$1379_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4148$1380_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4151$1381_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4154$1382_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4157$1383_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:416$136_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4160$1384_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4163$1385_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4166$1386_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4169$1387_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4172$1388_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4175$1389_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4178$1390_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4181$1391_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4184$1392_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4187$1393_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:419$137_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4190$1394_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4193$1395_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4196$1396_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4199$1397_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4202$1398_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4205$1399_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4208$1400_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4211$1401_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4214$1402_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4217$1403_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:422$138_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4220$1404_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4223$1405_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4226$1406_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4229$1407_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4232$1408_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4235$1409_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4238$1410_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4241$1411_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4244$1412_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4247$1413_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:425$139_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4250$1414_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4253$1415_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4256$1416_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4259$1417_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4262$1418_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4265$1419_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4268$1420_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4271$1421_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4274$1422_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4277$1423_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:428$140_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4280$1424_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4283$1425_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4286$1426_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4289$1427_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4292$1428_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4295$1429_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4298$1430_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4301$1431_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4304$1432_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4307$1433_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:431$141_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4310$1434_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4313$1435_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4316$1436_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4319$1437_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4322$1438_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4325$1439_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4328$1440_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4331$1441_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4334$1442_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4337$1443_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:434$142_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4340$1444_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4343$1445_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4346$1446_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4349$1447_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4352$1448_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4355$1449_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4358$1450_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4361$1451_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4364$1452_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4367$1453_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:437$143_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4370$1454_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4373$1455_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4376$1456_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4379$1457_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4382$1458_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4385$1459_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4388$1460_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4391$1461_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4394$1462_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4397$1463_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:440$144_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4400$1464_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4403$1465_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4406$1466_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4409$1467_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4412$1468_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4415$1469_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4418$1470_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4421$1471_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4424$1472_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4427$1473_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:443$145_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4430$1474_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4433$1475_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4436$1476_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4439$1477_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4442$1478_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4445$1479_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4448$1480_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4451$1481_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4454$1482_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4457$1483_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:446$146_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4460$1484_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4463$1485_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4466$1486_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4469$1487_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4472$1488_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4475$1489_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4478$1490_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4481$1491_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4484$1492_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4487$1493_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:449$147_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4490$1494_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4493$1495_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4496$1496_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4499$1497_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4502$1498_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4505$1499_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4508$1500_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4511$1501_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4514$1502_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4517$1503_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:452$148_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4520$1504_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4523$1505_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4526$1506_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4529$1507_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4532$1508_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4535$1509_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4538$1510_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4541$1511_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4544$1512_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4547$1513_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:455$149_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4550$1514_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4553$1515_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4556$1516_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4559$1517_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4562$1518_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4565$1519_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4568$1520_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4571$1521_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4574$1522_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4577$1523_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:458$150_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4580$1524_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4583$1525_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4586$1526_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4589$1527_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4592$1528_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4595$1529_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4598$1530_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4601$1531_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4604$1532_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4607$1533_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:461$151_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4610$1534_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4613$1535_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4616$1536_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4619$1537_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4622$1538_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4625$1539_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4628$1540_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4631$1541_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4634$1542_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4637$1543_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:464$152_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4640$1544_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4643$1545_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4646$1546_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4649$1547_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4652$1548_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4655$1549_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4658$1550_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4661$1551_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4664$1552_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4667$1553_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:467$153_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4670$1554_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4673$1555_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4676$1556_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4679$1557_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4682$1558_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4685$1559_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4688$1560_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4691$1561_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4694$1562_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4697$1563_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:470$154_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4700$1564_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4703$1565_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4706$1566_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4709$1567_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4712$1568_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4715$1569_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4718$1570_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4721$1571_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4724$1572_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4727$1573_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:473$155_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4730$1574_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4733$1575_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4736$1576_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4739$1577_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4742$1578_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4745$1579_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4748$1580_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4751$1581_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4754$1582_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4757$1583_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:476$156_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4760$1584_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4763$1585_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4766$1586_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4769$1587_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4772$1588_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4775$1589_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4778$1590_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4781$1591_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4784$1592_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4787$1593_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:479$157_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4790$1594_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4793$1595_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4796$1596_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4799$1597_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4802$1598_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4805$1599_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4808$1600_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4811$1601_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4814$1602_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4817$1603_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:482$158_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4820$1604_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4823$1605_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4826$1606_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4829$1607_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4832$1608_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4835$1609_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4838$1610_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4841$1611_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4844$1612_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4847$1613_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:485$159_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4850$1614_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4853$1615_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4856$1616_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4859$1617_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4862$1618_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4865$1619_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4868$1620_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4871$1621_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4874$1622_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4877$1623_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:488$160_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4880$1624_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4883$1625_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4886$1626_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4889$1627_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4892$1628_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4895$1629_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4898$1630_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4901$1631_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4904$1632_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4907$1633_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:491$161_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4910$1634_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4913$1635_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4916$1636_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4919$1637_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4922$1638_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4925$1639_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4928$1640_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4931$1641_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4934$1642_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4937$1643_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:494$162_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4940$1644_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4943$1645_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4946$1646_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4949$1647_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4952$1648_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4955$1649_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4958$1650_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4961$1651_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4964$1652_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4967$1653_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:497$163_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4970$1654_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4973$1655_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4976$1656_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4979$1657_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4982$1658_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4985$1659_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4988$1660_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4991$1661_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4994$1662_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:4997$1663_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:500$164_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5000$1664_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5003$1665_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5006$1666_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5009$1667_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5012$1668_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5015$1669_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5018$1670_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5021$1671_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5024$1672_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5027$1673_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:503$165_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5030$1674_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5033$1675_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5036$1676_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5039$1677_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5042$1678_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5045$1679_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5048$1680_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5051$1681_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5054$1682_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5057$1683_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:506$166_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5060$1684_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5063$1685_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5066$1686_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5069$1687_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5072$1688_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5075$1689_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5078$1690_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5081$1691_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5084$1692_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5087$1693_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:509$167_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5090$1694_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5093$1695_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5096$1696_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5099$1697_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5102$1698_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5105$1699_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5108$1700_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5111$1701_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5114$1702_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5117$1703_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:512$168_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5120$1704_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5123$1705_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5126$1706_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5129$1707_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5132$1708_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5135$1709_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5138$1710_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5141$1711_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5144$1712_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5147$1713_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:515$169_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5150$1714_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5153$1715_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5156$1716_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5159$1717_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5162$1718_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5165$1719_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5168$1720_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5171$1721_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5174$1722_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5177$1723_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:518$170_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5180$1724_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5183$1725_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5186$1726_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5189$1727_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5192$1728_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5195$1729_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5198$1730_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5201$1731_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5204$1732_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5207$1733_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:521$171_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5210$1734_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5213$1735_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5216$1736_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5219$1737_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5222$1738_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5225$1739_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5228$1740_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5231$1741_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5234$1742_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5237$1743_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:524$172_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5240$1744_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5243$1745_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5246$1746_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5249$1747_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5252$1748_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5255$1749_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5258$1750_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5261$1751_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5264$1752_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5267$1753_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:527$173_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5270$1754_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5273$1755_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5276$1756_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5279$1757_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5282$1758_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5285$1759_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5288$1760_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5291$1761_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5294$1762_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5297$1763_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:530$174_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5300$1764_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5303$1765_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5306$1766_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5309$1767_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5312$1768_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5315$1769_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5318$1770_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5321$1771_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5324$1772_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5327$1773_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:533$175_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5330$1774_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5333$1775_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5336$1776_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5339$1777_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5342$1778_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5345$1779_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5348$1780_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5351$1781_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5354$1782_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5357$1783_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:536$176_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5360$1784_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5363$1785_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5366$1786_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5369$1787_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5372$1788_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5375$1789_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5378$1790_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5381$1791_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5384$1792_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5387$1793_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:539$177_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5390$1794_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5393$1795_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5396$1796_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5399$1797_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5402$1798_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5405$1799_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5408$1800_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5411$1801_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5414$1802_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5417$1803_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:542$178_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5420$1804_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5423$1805_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5426$1806_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5429$1807_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5432$1808_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5435$1809_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5438$1810_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5441$1811_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5444$1812_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5447$1813_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:545$179_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5450$1814_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5453$1815_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5456$1816_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5459$1817_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5462$1818_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5465$1819_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5468$1820_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5471$1821_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5474$1822_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5477$1823_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:548$180_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5480$1824_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5483$1825_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5486$1826_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5489$1827_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5492$1828_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5495$1829_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5498$1830_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5501$1831_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5504$1832_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5507$1833_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:551$181_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5510$1834_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5513$1835_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5516$1836_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5519$1837_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5522$1838_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5525$1839_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5528$1840_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5531$1841_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5534$1842_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5537$1843_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:554$182_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5540$1844_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5543$1845_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5546$1846_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5549$1847_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5552$1848_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5555$1849_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5558$1850_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5561$1851_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5564$1852_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5567$1853_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:557$183_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5570$1854_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5573$1855_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5576$1856_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5579$1857_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5582$1858_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5585$1859_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5588$1860_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5591$1861_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5594$1862_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5597$1863_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:560$184_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5600$1864_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5603$1865_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5606$1866_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5609$1867_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5612$1868_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5615$1869_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5618$1870_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5621$1871_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5624$1872_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5627$1873_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:563$185_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5630$1874_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5633$1875_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5636$1876_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5639$1877_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5642$1878_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5645$1879_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5648$1880_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5651$1881_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5654$1882_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5657$1883_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:566$186_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5660$1884_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5663$1885_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5666$1886_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5669$1887_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5672$1888_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5675$1889_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5678$1890_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5681$1891_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5684$1892_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5687$1893_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:569$187_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5690$1894_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5693$1895_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5696$1896_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5699$1897_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5702$1898_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5705$1899_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5708$1900_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5711$1901_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5714$1902_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5717$1903_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:572$188_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5720$1904_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5723$1905_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5726$1906_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5729$1907_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5732$1908_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5735$1909_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5738$1910_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5741$1911_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5744$1912_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5747$1913_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:575$189_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5750$1914_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5753$1915_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5756$1916_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5759$1917_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5762$1918_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5765$1919_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5768$1920_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5771$1921_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5774$1922_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5777$1923_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:578$190_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5780$1924_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5783$1925_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5786$1926_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5789$1927_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5792$1928_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5795$1929_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5798$1930_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5801$1931_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5804$1932_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5807$1933_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:581$191_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5810$1934_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5813$1935_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5816$1936_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5819$1937_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5822$1938_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5825$1939_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5828$1940_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5831$1941_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5834$1942_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5837$1943_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:584$192_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5840$1944_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5843$1945_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5846$1946_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5849$1947_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5852$1948_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5855$1949_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5858$1950_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5861$1951_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5864$1952_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5867$1953_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:587$193_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5870$1954_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5873$1955_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5876$1956_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5879$1957_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5882$1958_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5885$1959_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5888$1960_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5891$1961_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5894$1962_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5897$1963_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:590$194_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5900$1964_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5903$1965_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5906$1966_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5909$1967_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5912$1968_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5915$1969_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5918$1970_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5921$1971_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5924$1972_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5927$1973_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:593$195_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5930$1974_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5933$1975_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5936$1976_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5939$1977_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5942$1978_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5945$1979_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5948$1980_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5951$1981_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5954$1982_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5957$1983_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:596$196_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5960$1984_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5963$1985_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5966$1986_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5969$1987_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5972$1988_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5975$1989_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5978$1990_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5981$1991_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5984$1992_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5987$1993_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:599$197_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5990$1994_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5993$1995_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5996$1996_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:5999$1997_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6002$1998_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6005$1999_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6008$2000_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6011$2001_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6014$2002_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6017$2003_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:602$198_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6020$2004_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6023$2005_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6026$2006_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6029$2007_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6032$2008_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6035$2009_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6038$2010_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6041$2011_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6044$2012_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6047$2013_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:605$199_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6050$2014_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6053$2015_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6056$2016_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6059$2017_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6062$2018_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6065$2019_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6068$2020_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6071$2021_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6074$2022_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6077$2023_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:608$200_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6080$2024_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6083$2025_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6086$2026_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6089$2027_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6092$2028_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6095$2029_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6098$2030_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6101$2031_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6104$2032_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6107$2033_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:611$201_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6110$2034_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6113$2035_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6116$2036_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6119$2037_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6122$2038_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6125$2039_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6128$2040_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6131$2041_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6134$2042_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6137$2043_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:614$202_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6140$2044_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6143$2045_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6146$2046_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6149$2047_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6152$2048_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6155$2049_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6158$2050_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6161$2051_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6164$2052_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6167$2053_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:617$203_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6170$2054_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6173$2055_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6176$2056_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6179$2057_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6182$2058_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6185$2059_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6188$2060_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6191$2061_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6194$2062_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6197$2063_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:620$204_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6200$2064_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6203$2065_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6206$2066_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6209$2067_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6212$2068_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6215$2069_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6218$2070_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6221$2071_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6224$2072_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6227$2073_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:623$205_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6230$2074_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6233$2075_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6236$2076_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6239$2077_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6242$2078_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6245$2079_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6248$2080_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6251$2081_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6254$2082_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6257$2083_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:626$206_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6260$2084_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6263$2085_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6266$2086_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6269$2087_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6272$2088_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6275$2089_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6278$2090_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6281$2091_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6284$2092_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6287$2093_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:629$207_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6290$2094_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6293$2095_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6296$2096_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6299$2097_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6302$2098_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6305$2099_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6308$2100_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6311$2101_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6314$2102_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6317$2103_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:632$208_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6320$2104_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6323$2105_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6326$2106_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6329$2107_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6332$2108_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6335$2109_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6338$2110_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6341$2111_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6344$2112_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6347$2113_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:635$209_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6350$2114_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6353$2115_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6356$2116_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6359$2117_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6362$2118_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6365$2119_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6368$2120_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6371$2121_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6374$2122_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6377$2123_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:638$210_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6380$2124_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6383$2125_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6386$2126_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6389$2127_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6392$2128_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6395$2129_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6398$2130_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6401$2131_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6404$2132_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6407$2133_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:641$211_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6410$2134_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6413$2135_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6416$2136_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6419$2137_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6422$2138_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6425$2139_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6428$2140_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6431$2141_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6434$2142_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6437$2143_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:644$212_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6440$2144_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6443$2145_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6446$2146_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6449$2147_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6452$2148_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6455$2149_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6458$2150_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6461$2151_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6464$2152_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6467$2153_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:647$213_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6470$2154_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6473$2155_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6476$2156_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6479$2157_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6482$2158_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6485$2159_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6488$2160_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6491$2161_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6494$2162_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6497$2163_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:650$214_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6500$2164_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6503$2165_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6506$2166_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6509$2167_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6512$2168_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6515$2169_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6518$2170_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6521$2171_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6524$2172_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6527$2173_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:653$215_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6530$2174_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6533$2175_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6536$2176_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6539$2177_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6542$2178_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6545$2179_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6548$2180_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6551$2181_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6554$2182_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6557$2183_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:656$216_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6560$2184_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6563$2185_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6566$2186_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6569$2187_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6572$2188_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6575$2189_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6578$2190_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6581$2191_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6584$2192_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6587$2193_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:659$217_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6590$2194_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6593$2195_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6596$2196_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6599$2197_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6602$2198_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6605$2199_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6608$2200_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6611$2201_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6614$2202_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6617$2203_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:662$218_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6620$2204_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6623$2205_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6626$2206_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6629$2207_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6632$2208_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6635$2209_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6638$2210_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6641$2211_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6644$2212_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6647$2213_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:665$219_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6650$2214_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6653$2215_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6656$2216_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6659$2217_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6662$2218_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6665$2219_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6668$2220_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6671$2221_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6674$2222_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6677$2223_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:668$220_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6680$2224_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6683$2225_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6686$2226_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6689$2227_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6692$2228_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6695$2229_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6698$2230_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6701$2231_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6704$2232_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6707$2233_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:671$221_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6710$2234_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6713$2235_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6716$2236_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6719$2237_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6722$2238_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6725$2239_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6728$2240_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6731$2241_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6734$2242_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6737$2243_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:674$222_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6740$2244_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6743$2245_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6746$2246_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6749$2247_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6752$2248_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6755$2249_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6758$2250_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6761$2251_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6764$2252_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6767$2253_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:677$223_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6770$2254_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6773$2255_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6776$2256_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6779$2257_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6782$2258_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6785$2259_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6788$2260_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6791$2261_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6794$2262_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6797$2263_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:680$224_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6800$2264_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6803$2265_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6806$2266_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6809$2267_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6812$2268_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6815$2269_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6818$2270_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6821$2271_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6824$2272_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6827$2273_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:683$225_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6830$2274_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6833$2275_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6836$2276_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6839$2277_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6842$2278_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6845$2279_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6848$2280_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6851$2281_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6854$2282_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6857$2283_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:686$226_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6860$2284_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6863$2285_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6866$2286_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6869$2287_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6872$2288_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6875$2289_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6878$2290_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6881$2291_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6884$2292_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6887$2293_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:689$227_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6890$2294_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6893$2295_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6896$2296_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6899$2297_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6902$2298_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6905$2299_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6908$2300_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6911$2301_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6914$2302_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6917$2303_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:692$228_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6920$2304_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6923$2305_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6926$2306_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6929$2307_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6932$2308_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6935$2309_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6938$2310_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6941$2311_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6944$2312_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6947$2313_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:695$229_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6950$2314_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6953$2315_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6956$2316_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6959$2317_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6962$2318_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6965$2319_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6968$2320_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6971$2321_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6974$2322_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6977$2323_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:698$230_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6980$2324_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6983$2325_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6986$2326_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6989$2327_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6992$2328_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6995$2329_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:6998$2330_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7001$2331_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7004$2332_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7007$2333_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:701$231_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7010$2334_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7013$2335_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7016$2336_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7019$2337_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7022$2338_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7025$2339_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7028$2340_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7031$2341_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7034$2342_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7037$2343_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:704$232_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7040$2344_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7043$2345_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7046$2346_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7049$2347_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7052$2348_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7055$2349_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7058$2350_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7061$2351_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7064$2352_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7067$2353_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:707$233_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7070$2354_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7073$2355_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7076$2356_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7079$2357_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7082$2358_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7085$2359_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7088$2360_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7091$2361_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7094$2362_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7097$2363_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:710$234_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7100$2364_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7103$2365_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7106$2366_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7109$2367_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7112$2368_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7115$2369_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7118$2370_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7121$2371_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7124$2372_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7127$2373_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:713$235_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7130$2374_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7133$2375_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7136$2376_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7139$2377_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7142$2378_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7145$2379_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7148$2380_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7151$2381_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7154$2382_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7157$2383_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:716$236_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7160$2384_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7163$2385_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7166$2386_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7169$2387_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7172$2388_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7175$2389_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7178$2390_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7181$2391_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7184$2392_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7187$2393_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:719$237_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7190$2394_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7193$2395_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7196$2396_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7199$2397_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7202$2398_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7205$2399_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7208$2400_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7211$2401_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7214$2402_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7217$2403_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:722$238_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7220$2404_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7223$2405_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7226$2406_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7229$2407_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7232$2408_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7235$2409_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7238$2410_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7241$2411_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7244$2412_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7247$2413_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:725$239_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7250$2414_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7253$2415_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7256$2416_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7259$2417_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7262$2418_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7265$2419_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7268$2420_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7271$2421_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7274$2422_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7277$2423_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:728$240_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7280$2424_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7283$2425_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7286$2426_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7289$2427_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7292$2428_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7295$2429_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7298$2430_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7301$2431_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7304$2432_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7307$2433_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:731$241_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7310$2434_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7313$2435_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7316$2436_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7319$2437_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7322$2438_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7325$2439_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7328$2440_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7331$2441_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7334$2442_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7337$2443_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:734$242_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7340$2444_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7343$2445_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7346$2446_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7349$2447_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7352$2448_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7355$2449_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7358$2450_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7361$2451_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7364$2452_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7367$2453_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:737$243_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7370$2454_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7373$2455_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7376$2456_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7379$2457_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7382$2458_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7385$2459_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7388$2460_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7391$2461_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7394$2462_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7397$2463_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:740$244_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7400$2464_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7403$2465_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7406$2466_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7409$2467_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7412$2468_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7415$2469_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7418$2470_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7421$2471_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7424$2472_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7427$2473_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:743$245_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7430$2474_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7433$2475_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7436$2476_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7439$2477_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7442$2478_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7445$2479_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7448$2480_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7451$2481_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7454$2482_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7457$2483_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:746$246_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7460$2484_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7463$2485_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7466$2486_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7469$2487_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7472$2488_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7475$2489_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7478$2490_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7481$2491_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7484$2492_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7487$2493_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:749$247_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7490$2494_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7493$2495_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7496$2496_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7499$2497_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7502$2498_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7505$2499_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7508$2500_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7511$2501_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7514$2502_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7517$2503_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:752$248_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7520$2504_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7523$2505_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7526$2506_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7529$2507_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7532$2508_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7535$2509_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7538$2510_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7541$2511_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7544$2512_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7547$2513_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:755$249_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7550$2514_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7553$2515_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7556$2516_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7559$2517_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7562$2518_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7565$2519_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7568$2520_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7571$2521_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7574$2522_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7577$2523_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:758$250_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7580$2524_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7583$2525_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7586$2526_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7589$2527_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7592$2528_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7595$2529_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7598$2530_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7601$2531_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7604$2532_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7607$2533_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:761$251_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7610$2534_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7613$2535_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7616$2536_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7619$2537_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7622$2538_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7625$2539_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7628$2540_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7631$2541_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7634$2542_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7637$2543_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:764$252_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7640$2544_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7643$2545_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7646$2546_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7649$2547_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7652$2548_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7655$2549_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7658$2550_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7661$2551_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7664$2552_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7667$2553_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:767$253_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7670$2554_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7673$2555_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7676$2556_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7679$2557_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7682$2558_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7685$2559_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7688$2560_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7691$2561_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7694$2562_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7697$2563_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:770$254_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7700$2564_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7703$2565_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7706$2566_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7709$2567_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7712$2568_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7715$2569_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7718$2570_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7721$2571_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7724$2572_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7727$2573_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:773$255_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7730$2574_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7733$2575_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7736$2576_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7739$2577_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7742$2578_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7745$2579_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7748$2580_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7751$2581_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7754$2582_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7757$2583_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:776$256_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7760$2584_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7763$2585_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7766$2586_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7769$2587_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7772$2588_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7775$2589_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7778$2590_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7781$2591_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7784$2592_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7787$2593_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:779$257_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7790$2594_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7793$2595_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7796$2596_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7799$2597_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7802$2598_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7805$2599_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7808$2600_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7811$2601_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7814$2602_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7817$2603_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:782$258_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7820$2604_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7823$2605_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7826$2606_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7829$2607_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7832$2608_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7835$2609_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7838$2610_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7841$2611_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7844$2612_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7847$2613_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:785$259_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7850$2614_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7853$2615_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7856$2616_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7859$2617_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7862$2618_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7865$2619_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7868$2620_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7871$2621_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7874$2622_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7877$2623_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:788$260_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7880$2624_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7883$2625_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7886$2626_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7889$2627_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7892$2628_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7895$2629_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7898$2630_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7901$2631_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7904$2632_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7907$2633_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:791$261_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7910$2634_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7913$2635_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7916$2636_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7919$2637_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7922$2638_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7925$2639_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7928$2640_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7931$2641_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7934$2642_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7937$2643_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:794$262_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7940$2644_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7943$2645_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7946$2646_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7949$2647_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7952$2648_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7955$2649_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7958$2650_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7961$2651_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7964$2652_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7967$2653_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:797$263_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7970$2654_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7973$2655_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7976$2656_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7979$2657_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7982$2658_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7985$2659_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7988$2660_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7991$2661_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7994$2662_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:7997$2663_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:800$264_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8000$2664_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8003$2665_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8006$2666_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8009$2667_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8012$2668_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8015$2669_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8018$2670_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8021$2671_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8024$2672_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8027$2673_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:803$265_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8030$2674_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8033$2675_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8036$2676_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8039$2677_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8042$2678_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8045$2679_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8048$2680_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8051$2681_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8054$2682_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8057$2683_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:806$266_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8060$2684_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8063$2685_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8066$2686_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8069$2687_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8072$2688_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8075$2689_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8078$2690_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8081$2691_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8084$2692_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8087$2693_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:809$267_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8090$2694_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8093$2695_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8096$2696_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8099$2697_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8102$2698_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8105$2699_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8108$2700_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8111$2701_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8114$2702_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8117$2703_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:812$268_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8120$2704_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8123$2705_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8126$2706_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8129$2707_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8132$2708_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8135$2709_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8138$2710_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8141$2711_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8144$2712_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8147$2713_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:815$269_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8150$2714_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8153$2715_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8156$2716_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8159$2717_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8162$2718_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8165$2719_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8168$2720_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8171$2721_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8174$2722_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8177$2723_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:818$270_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8180$2724_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8183$2725_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8186$2726_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8189$2727_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8192$2728_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8195$2729_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8198$2730_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8201$2731_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8204$2732_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8207$2733_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:821$271_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8210$2734_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8213$2735_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8216$2736_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8219$2737_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8222$2738_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8225$2739_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8228$2740_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8231$2741_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8234$2742_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8237$2743_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:824$272_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8240$2744_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8243$2745_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8246$2746_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8249$2747_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8252$2748_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8255$2749_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8258$2750_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8261$2751_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8264$2752_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8267$2753_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:827$273_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8270$2754_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8273$2755_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8276$2756_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8279$2757_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8282$2758_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8285$2759_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8288$2760_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8291$2761_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8294$2762_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8297$2763_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:830$274_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8300$2764_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8303$2765_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8306$2766_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8309$2767_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8312$2768_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8315$2769_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8318$2770_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8321$2771_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8324$2772_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8327$2773_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:833$275_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8330$2774_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8333$2775_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8336$2776_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8339$2777_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8342$2778_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8345$2779_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8348$2780_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8351$2781_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8354$2782_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8357$2783_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:836$276_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8360$2784_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8363$2785_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8366$2786_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8369$2787_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8372$2788_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8375$2789_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8378$2790_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8381$2791_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8384$2792_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8387$2793_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:839$277_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8390$2794_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8393$2795_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8396$2796_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8399$2797_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8402$2798_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8405$2799_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8408$2800_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8411$2801_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8414$2802_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8417$2803_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:842$278_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8420$2804_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8423$2805_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8426$2806_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8429$2807_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8432$2808_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8435$2809_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8438$2810_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8441$2811_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8444$2812_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8447$2813_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:845$279_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8450$2814_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8453$2815_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8456$2816_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8459$2817_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8462$2818_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8465$2819_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8468$2820_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8471$2821_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8474$2822_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8477$2823_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:848$280_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8480$2824_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8483$2825_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8486$2826_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8489$2827_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8492$2828_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8495$2829_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8498$2830_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8501$2831_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8504$2832_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8507$2833_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:851$281_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8510$2834_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8513$2835_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8516$2836_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8519$2837_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8522$2838_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8525$2839_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8528$2840_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8531$2841_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8534$2842_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8537$2843_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:854$282_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8540$2844_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8543$2845_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8546$2846_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8549$2847_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8552$2848_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8555$2849_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8558$2850_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8561$2851_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8564$2852_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8567$2853_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:857$283_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8570$2854_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8573$2855_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8576$2856_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8579$2857_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8582$2858_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8585$2859_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8588$2860_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8591$2861_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8594$2862_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8597$2863_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:860$284_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8600$2864_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8603$2865_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8606$2866_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8609$2867_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8612$2868_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8615$2869_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8618$2870_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8621$2871_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8624$2872_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8627$2873_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:863$285_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8630$2874_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8633$2875_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8636$2876_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8639$2877_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8642$2878_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8645$2879_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8648$2880_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8651$2881_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8654$2882_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8657$2883_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:866$286_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8660$2884_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8663$2885_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8666$2886_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8669$2887_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8672$2888_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8675$2889_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8678$2890_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8681$2891_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8684$2892_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8687$2893_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:869$287_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8690$2894_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8693$2895_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8696$2896_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8699$2897_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8702$2898_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8705$2899_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8708$2900_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8711$2901_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8714$2902_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8717$2903_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:872$288_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8720$2904_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8723$2905_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8726$2906_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8729$2907_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8732$2908_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8735$2909_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8738$2910_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8741$2911_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8744$2912_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8747$2913_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:875$289_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8750$2914_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8753$2915_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8756$2916_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8759$2917_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8762$2918_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8765$2919_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8768$2920_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8771$2921_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8774$2922_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8777$2923_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:878$290_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8780$2924_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8783$2925_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8786$2926_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8789$2927_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8792$2928_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8795$2929_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8798$2930_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8801$2931_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8804$2932_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8807$2933_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:881$291_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8810$2934_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8813$2935_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8816$2936_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8819$2937_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8822$2938_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8825$2939_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8828$2940_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8831$2941_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8834$2942_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8837$2943_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:884$292_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8840$2944_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8843$2945_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8846$2946_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8849$2947_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8852$2948_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8855$2949_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8858$2950_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8861$2951_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8864$2952_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8867$2953_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:887$293_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8870$2954_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8873$2955_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8876$2956_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8879$2957_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8882$2958_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8885$2959_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8888$2960_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8891$2961_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8894$2962_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8897$2963_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:890$294_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8900$2964_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8903$2965_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8906$2966_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8909$2967_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8912$2968_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8915$2969_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8918$2970_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8921$2971_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8924$2972_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8927$2973_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:893$295_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8930$2974_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8933$2975_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8936$2976_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8939$2977_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8942$2978_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8945$2979_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8948$2980_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8951$2981_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8954$2982_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8957$2983_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:896$296_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8960$2984_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8963$2985_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8966$2986_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8969$2987_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8972$2988_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8975$2989_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8978$2990_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8981$2991_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8984$2992_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8987$2993_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:899$297_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8990$2994_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8993$2995_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8996$2996_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:8999$2997_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9002$2998_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9005$2999_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9008$3000_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9011$3001_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9014$3002_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9017$3003_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:902$298_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9020$3004_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9023$3005_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9026$3006_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9029$3007_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9032$3008_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9035$3009_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9038$3010_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9041$3011_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9044$3012_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9047$3013_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:905$299_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9050$3014_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9053$3015_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9056$3016_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9059$3017_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9062$3018_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9065$3019_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9068$3020_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9071$3021_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9074$3022_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9077$3023_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:908$300_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9080$3024_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9083$3025_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9086$3026_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9089$3027_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9092$3028_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9095$3029_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9098$3030_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9101$3031_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9104$3032_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9107$3033_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:911$301_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9110$3034_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9113$3035_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9116$3036_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9119$3037_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9122$3038_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9125$3039_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9128$3040_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9131$3041_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9134$3042_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9137$3043_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:914$302_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9140$3044_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9143$3045_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9146$3046_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9149$3047_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9152$3048_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9155$3049_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9158$3050_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9161$3051_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9164$3052_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9167$3053_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:917$303_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9170$3054_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9173$3055_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9176$3056_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9179$3057_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9182$3058_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9185$3059_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9188$3060_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9191$3061_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9194$3062_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9197$3063_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:920$304_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9200$3064_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9203$3065_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9206$3066_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9209$3067_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9212$3068_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9215$3069_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9218$3070_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9221$3071_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9224$3072_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9227$3073_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:923$305_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9230$3074_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9233$3075_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9236$3076_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9239$3077_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9242$3078_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9245$3079_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9248$3080_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9251$3081_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9254$3082_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9257$3083_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:926$306_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9260$3084_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9263$3085_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9266$3086_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9269$3087_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9272$3088_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9275$3089_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9278$3090_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9281$3091_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9284$3092_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9287$3093_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:929$307_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9290$3094_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9293$3095_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9296$3096_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9299$3097_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9302$3098_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9305$3099_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9308$3100_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9311$3101_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9314$3102_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9317$3103_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:932$308_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9320$3104_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9323$3105_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9326$3106_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9329$3107_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9332$3108_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9335$3109_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9338$3110_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9341$3111_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9344$3112_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9347$3113_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:935$309_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9350$3114_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9353$3115_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9356$3116_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9359$3117_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9362$3118_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9365$3119_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9368$3120_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9371$3121_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9374$3122_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9377$3123_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:938$310_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9380$3124_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9383$3125_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9386$3126_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9389$3127_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9392$3128_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9395$3129_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9398$3130_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9401$3131_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9404$3132_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9407$3133_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:941$311_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9410$3134_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9413$3135_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9416$3136_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9419$3137_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9422$3138_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9425$3139_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9428$3140_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9431$3141_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9434$3142_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9437$3143_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:944$312_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9440$3144_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9443$3145_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9446$3146_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9449$3147_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9452$3148_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9455$3149_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9458$3150_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9461$3151_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9464$3152_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9467$3153_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:947$313_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9470$3154_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9473$3155_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9476$3156_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9479$3157_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9482$3158_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9485$3159_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9488$3160_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9491$3161_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9494$3162_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9497$3163_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:950$314_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9500$3164_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9503$3165_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9506$3166_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9509$3167_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9512$3168_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9515$3169_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9518$3170_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9521$3171_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9524$3172_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9527$3173_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:953$315_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9530$3174_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9533$3175_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9536$3176_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9539$3177_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9542$3178_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9545$3179_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9548$3180_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9551$3181_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9554$3182_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9557$3183_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:956$316_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9560$3184_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9563$3185_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9566$3186_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9569$3187_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9572$3188_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9575$3189_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9578$3190_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9581$3191_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9584$3192_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9587$3193_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:959$317_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9590$3194_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9593$3195_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9596$3196_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9599$3197_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9602$3198_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9605$3199_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9608$3200_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9611$3201_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9614$3202_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9617$3203_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:962$318_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9620$3204_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9623$3205_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9626$3206_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9629$3207_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9632$3208_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9635$3209_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9638$3210_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9641$3211_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9644$3212_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9647$3213_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:965$319_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9650$3214_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9653$3215_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9656$3216_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9659$3217_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9662$3218_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9665$3219_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9668$3220_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9671$3221_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9674$3222_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9677$3223_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:968$320_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9680$3224_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9683$3225_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9686$3226_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9689$3227_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9692$3228_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9695$3229_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9698$3230_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9701$3231_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9704$3232_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9707$3233_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:971$321_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9710$3234_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9713$3235_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9716$3236_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9719$3237_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9722$3238_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9725$3239_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9728$3240_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9731$3241_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9734$3242_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9737$3243_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:974$322_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9740$3244_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9743$3245_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9746$3246_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9749$3247_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9752$3248_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9755$3249_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9758$3250_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9761$3251_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9764$3252_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9767$3253_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:977$323_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9770$3254_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9773$3255_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9776$3256_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9779$3257_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9782$3258_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9785$3259_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9788$3260_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9791$3261_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9794$3262_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9797$3263_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:980$324_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9800$3264_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9803$3265_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9806$3266_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9809$3267_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9812$3268_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9815$3269_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9818$3270_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9821$3271_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9824$3272_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9827$3273_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:983$325_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9830$3274_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9833$3275_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9836$3276_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9839$3277_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9842$3278_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9845$3279_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9848$3280_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9851$3281_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9854$3282_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9857$3283_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:986$326_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9860$3284_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9863$3285_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9866$3286_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9869$3287_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9872$3288_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9875$3289_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9878$3290_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9881$3291_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9884$3292_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9887$3293_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:989$327_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9890$3294_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9893$3295_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9896$3296_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9899$3297_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9902$3298_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9905$3299_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9908$3300_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9911$3301_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9914$3302_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9917$3303_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:992$328_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9920$3304_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9923$3305_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9926$3306_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9929$3307_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9932$3308_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9935$3309_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9938$3310_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9941$3311_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9944$3312_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9947$3313_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:995$329_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9950$3314_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9953$3315_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9956$3316_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9959$3317_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9962$3318_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9965$3319_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9968$3320_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9971$3321_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9974$3322_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9977$3323_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:998$330_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9980$3324_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9983$3325_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9986$3326_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9989$3327_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9992$3328_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9995$3329_CHECK  = 1'b0;
    // UUT.tracker.$formal$SignalTracker.\sv:9998$3330_CHECK  = 1'b0;
    UUT._mem[20'b00000000000000000000] = 64'b0000000101000010001010000011001100000010011100100100101011100011;
    UUT._mem[20'b00000000000001000000] = 64'b0000000101001010001010000011001111111111101000001110101000010011;
    UUT._mem[20'b00000000000001000001] = 64'b0001000000100000000000000111001100000000000000000000000001110011;
    UUT._mem[20'b00000000000001000010] = 64'b0000000101000010001010000011001100000010011100100100101011100011;
    UUT.dut.core.dpath.regFile.regs[5'b00000] = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.regFile.regs[5'b11010] = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.regFile.regs[5'b00001] = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.regFile.regs[5'b10100] = 32'b00000000000000000000000000000000;
    UUT.dut.core.dpath.regFile.regs[5'b00010] = 32'b00000000000000000000000000000000;
    UUT.dut.dcache.dataMem_0_0[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_0_1[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_0_2[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_0_3[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_1_0[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_1_1[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_1_2[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_1_3[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_2_0[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_2_1[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_2_2[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_2_3[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_3_0[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_3_1[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_3_2[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.dataMem_3_3[8'b00000000] = 8'b00000000;
    UUT.dut.dcache.metaMem_tag[8'b00000000] = 20'b00000000000000000000;
    UUT.dut.icache.dataMem_0_0[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_0_0[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_0_0[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_0_1[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_0_1[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_0_1[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_0_2[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_0_2[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_0_2[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_0_3[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_0_3[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_0_3[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_1_0[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_1_0[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_1_0[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_1_1[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_1_1[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_1_1[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_1_2[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_1_2[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_1_2[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_1_3[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_1_3[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_1_3[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_2_0[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_2_0[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_2_0[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_2_1[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_2_1[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_2_1[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_2_2[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_2_2[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_2_2[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_2_3[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_2_3[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_2_3[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_3_0[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_3_0[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_3_0[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_3_1[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_3_1[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_3_1[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_3_2[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_3_2[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_3_2[8'b00100001] = 8'b00000000;
    UUT.dut.icache.dataMem_3_3[8'b00000000] = 8'b00000000;
    UUT.dut.icache.dataMem_3_3[8'b00100000] = 8'b00000000;
    UUT.dut.icache.dataMem_3_3[8'b00100001] = 8'b00000000;
    UUT.dut.icache.metaMem_tag[8'b00000000] = 20'b00000000000000000000;
    UUT.dut.icache.metaMem_tag[8'b00100000] = 20'b00000000000000000000;
    UUT.dut.icache.metaMem_tag[8'b00100001] = 20'b00000000000000000000;

    // state 0
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
    end

    // state 2
    if (cycle == 1) begin
    end

    // state 3
    if (cycle == 2) begin
    end

    // state 4
    if (cycle == 3) begin
    end

    // state 5
    if (cycle == 4) begin
    end

    // state 6
    if (cycle == 5) begin
    end

    // state 7
    if (cycle == 6) begin
    end

    // state 8
    if (cycle == 7) begin
    end

    // state 9
    if (cycle == 8) begin
    end

    // state 10
    if (cycle == 9) begin
    end

    genclock <= cycle < 10;
    cycle <= cycle + 1;
  end
endmodule
