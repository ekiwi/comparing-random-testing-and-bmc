module SignalTracker(
  input clock,
  input reset,
  input dut__core__dpath__csr___io_out_T_29_0,
  input dut__core__dpath__csr___T_0,
  input dut__core__dpath__csr__isInstRet_0,
  input dut__core__dpath__csr___T_10_0,
  input dut__core__dpath__csr___T_7_0,
  input dut__core__dpath__csr___io_out_T_33_0,
  input dut__core__dpath__csr___T_23_0,
  input dut__core__dpath__csr___io_out_T_25_0,
  input dut__core__dpath__csr___T_6_0,
  input dut__core__dpath__csr___io_out_T_31_0,
  input dut__core__dpath__csr___wdata_T_3_0,
  input dut__core__dpath__csr__privInst_0,
  input dut__core__dpath__csr___T_16_0,
  input dut__core__dpath__csr__isEret_0,
  input dut__core__dpath__csr___io_out_T_41_0,
  input dut__core__dpath__csr___io_out_T_1_0,
  input dut__core__dpath__csr___io_out_T_53_0,
  input dut__core__dpath__csr__iaddrInvalid_0,
  input dut__core__dpath__csr___io_out_T_27_0,
  input dut__core__dpath__csr___io_out_T_43_0,
  input dut__core__dpath__csr___T_1_0,
  input dut__core__dpath__csr___io_out_T_35_0,
  input dut__core__dpath__csr___T_3_0,
  input dut__core__dpath__csr___T_18_0,
  input dut__core__dpath__csr__privValid_0,
  input dut__core__dpath__csr___io_expt_T_6_0,
  input dut__core__dpath__csr___isInstRet_T_0,
  input dut__core__dpath__csr___io_out_T_3_0,
  input dut__core__dpath__csr___io_out_T_7_0,
  input dut__core__dpath__csr__io_expt_0,
  input dut__core__dpath__csr___T_24_0,
  input dut__core__dpath__csr___wen_T_0,
  input dut__core__dpath__csr___T_21_0,
  input dut__core__dpath__csr__wen_0,
  input dut__core__dpath__csr___T_13_0,
  input dut__core__dpath__csr___T_8_0,
  input dut__core__dpath__csr___io_out_T_47_0,
  input dut__core__dpath__csr___io_out_T_19_0,
  input dut__core__dpath__csr___T_12_0,
  input dut__core__dpath__csr___io_out_T_9_0,
  input dut__core__dpath__csr___csrRO_T_4_0,
  input dut__core__dpath__csr___io_out_T_5_0,
  input dut__core__dpath__csr___isEcall_T_1_0,
  input dut__core__dpath__csr___wdata_T_5_0,
  input dut__core__dpath__csr___laddrInvalid_T_6_0,
  input dut__core__dpath__csr___T_17_0,
  input dut__core__dpath__csr___laddrInvalid_T_8_0,
  input dut__core__dpath__csr___io_out_T_45_0,
  input dut__core__dpath__csr___io_out_T_17_0,
  input dut__core__dpath__csr___io_out_T_13_0,
  input dut__core__dpath__csr___io_out_T_11_0,
  input dut__core__dpath__csr___T_20_0,
  input dut__core__dpath__csr___T_14_0,
  input dut__core__dpath__csr___io_out_T_55_0,
  input dut__core__dpath__csr___io_out_T_39_0,
  input dut__core__dpath__csr___io_out_T_51_0,
  input dut__core__dpath__csr__laddrInvalid_0,
  input dut__core__dpath__csr___io_out_T_23_0,
  input dut__core__dpath__csr___isInstRet_T_1_0,
  input dut__core__dpath__csr___io_expt_T_5_0,
  input dut__core__dpath__csr___isEcall_T_4_0,
  input dut__core__dpath__csr___csrRO_T_2_0,
  input dut__core__dpath__csr___saddrInvalid_T_3_0,
  input dut__core__dpath__csr__isEcall_0,
  input dut__core__dpath__csr__isEbreak_0,
  input dut__core__dpath__csr___io_out_T_49_0,
  input dut__core__dpath__csr___T_11_0,
  input dut__core__dpath__csr___wdata_T_7_0,
  input dut__core__dpath__csr___isInstRet_T_5_0,
  input dut__core__dpath__csr___io_out_T_37_0,
  input dut__core__dpath__csr___saddrInvalid_T_5_0,
  input dut__core__dpath__csr___T_22_0,
  input dut__core__dpath__csr___io_out_T_57_0,
  input dut__core__dpath__csr___laddrInvalid_T_4_0,
  input dut__core__dpath__csr___T_9_0,
  input dut__core__dpath__csr___T_15_0,
  input dut__core__dpath__csr__saddrInvalid_0,
  input dut__core__dpath__csr___T_19_0,
  input dut__core__dpath__csr___io_out_T_21_0,
  input dut__core__dpath__csr___io_out_T_15_0,
  input dut__core__dpath__regFile___T_1_0,
  input dut__core__dpath__regFile___io_rdata2_T_0,
  input dut__core__dpath__regFile___io_rdata1_T_0,
  input dut__core__dpath__alu___out_T_1_0,
  input dut__core__dpath__alu___cmp_T_4_0,
  input dut__core__dpath__alu___out_T_0,
  input dut__core__dpath__alu___out_T_10_0,
  input dut__core__dpath__alu___out_T_12_0,
  input dut__core__dpath__alu___shin_T_0,
  input dut__core__dpath__alu___out_T_9_0,
  input dut__core__dpath__alu___out_T_4_0,
  input dut__core__dpath__alu___out_T_3_0,
  input dut__core__dpath__alu___out_T_14_0,
  input dut__core__dpath__alu___out_T_6_0,
  input dut__core__dpath__alu___out_T_7_0,
  input dut__core__dpath__alu___out_T_8_0,
  input dut__core__dpath__alu___cmp_T_2_0,
  input dut__core__dpath__alu___sum_T_0,
  input dut__core__dpath__alu___out_T_5_0,
  input dut__core__dpath__alu___out_T_2_0,
  input dut__core__dpath__alu___out_T_16_0,
  input dut__core__dpath__immGen___io_out_T_2_0,
  input dut__core__dpath__immGen___io_out_T_4_0,
  input dut__core__dpath__immGen___io_out_T_6_0,
  input dut__core__dpath__immGen___io_out_T_12_0,
  input dut__core__dpath__immGen___io_out_T_8_0,
  input dut__core__dpath__immGen___io_out_T_10_0,
  input dut__core__dpath__brCond__isSameSign_0,
  input dut__core__dpath__brCond__eq_0,
  input dut__core__dpath__brCond___io_taken_T_5_0,
  input dut__core__dpath__brCond___io_taken_T_0,
  input dut__core__dpath__brCond___io_taken_T_11_0,
  input dut__core__dpath__brCond___io_taken_T_8_0,
  input dut__core__dpath__brCond___io_taken_T_14_0,
  input dut__core__dpath__brCond___io_taken_T_2_0,
  input dut__core__dpath__brCond__geu_0,
  input dut__core__dpath__brCond__ge_0,
  input dut__core__dpath___io_dcache_req_bits_mask_T_7_0,
  input dut__core__dpath___npc_T_2_0,
  input dut__core__dpath___inst_T_2_0,
  input dut__core__dpath___rs1_T_0,
  input dut__core__dpath___T_6_0,
  input dut__core__dpath__io_ctrl_A_sel_0,
  input dut__core__dpath___npc_T_5_0,
  input dut__core__dpath___io_icache_req_valid_T_0,
  input dut__core__dpath__io_ctrl_B_sel_0,
  input dut__core__dpath___regWrite_T_9_0,
  input dut__core__dpath___stall_T_1_0,
  input dut__core__dpath__csr__io_expt,
  input dut__core__dpath___regWrite_T_7_0,
  input dut__core__dpath___stall_T_0,
  input dut__core__dpath___rs1hazard_T_2_0,
  input dut__core__dpath___load_T_13_0,
  input dut__core__dpath___load_T_11_0,
  input dut__core__dpath___rs1_T_1_0,
  input dut__core__dpath__stall_0,
  input dut__core__dpath___io_dcache_req_bits_mask_T_9_0,
  input dut__core__dpath___load_T_15_0,
  input dut__core__dpath___io_dcache_req_bits_mask_T_5_0,
  input dut__core__dpath___rs2hazard_T_2_0,
  input dut__core__dpath___csr_in_T_0,
  input dut__core__dpath___npc_T_0,
  input dut__core__dpath___regWrite_T_5_0,
  input dut__core__dpath___npc_T_1_0,
  input dut__core__dpath___rs2_T_1_0,
  input dut__core__dpath___load_T_9_0,
  input dut__core__dpath___T_4_0,
  input dut__core__dpath___T_7_0,
  input dut__core__ctrl___ctrlSignals_T_31_0,
  input dut__core__ctrl___ctrlSignals_T_93_0,
  input dut__core__ctrl___ctrlSignals_T_87_0,
  input dut__core__ctrl___ctrlSignals_T_81_0,
  input dut__core__ctrl___ctrlSignals_T_15_0,
  input dut__core__ctrl___ctrlSignals_T_49_0,
  input dut__core__ctrl___ctrlSignals_T_5_0,
  input dut__core__ctrl___ctrlSignals_T_41_0,
  input dut__core__ctrl___ctrlSignals_T_11_0,
  input dut__core__ctrl___ctrlSignals_T_19_0,
  input dut__core__ctrl___ctrlSignals_T_95_0,
  input dut__core__ctrl___ctrlSignals_T_21_0,
  input dut__core__ctrl___ctrlSignals_T_47_0,
  input dut__core__ctrl___ctrlSignals_T_35_0,
  input dut__core__ctrl___ctrlSignals_T_75_0,
  input dut__core__ctrl___ctrlSignals_T_25_0,
  input dut__core__ctrl___ctrlSignals_T_55_0,
  input dut__core__ctrl___ctrlSignals_T_71_0,
  input dut__core__ctrl___ctrlSignals_T_27_0,
  input dut__core__ctrl___ctrlSignals_T_59_0,
  input dut__core__ctrl___ctrlSignals_T_29_0,
  input dut__core__ctrl___ctrlSignals_T_39_0,
  input dut__core__ctrl___ctrlSignals_T_1_0,
  input dut__core__ctrl___ctrlSignals_T_63_0,
  input dut__core__ctrl___ctrlSignals_T_97_0,
  input dut__core__ctrl___ctrlSignals_T_23_0,
  input dut__core__ctrl___ctrlSignals_T_65_0,
  input dut__core__ctrl___ctrlSignals_T_89_0,
  input dut__core__ctrl___ctrlSignals_T_51_0,
  input dut__core__ctrl___ctrlSignals_T_83_0,
  input dut__core__ctrl___ctrlSignals_T_77_0,
  input dut__core__ctrl___ctrlSignals_T_85_0,
  input dut__core__ctrl___ctrlSignals_T_37_0,
  input dut__core__ctrl___ctrlSignals_T_67_0,
  input dut__core__ctrl___ctrlSignals_T_91_0,
  input dut__core__ctrl___ctrlSignals_T_43_0,
  input dut__core__ctrl___ctrlSignals_T_17_0,
  input dut__core__ctrl___ctrlSignals_T_9_0,
  input dut__core__ctrl___ctrlSignals_T_79_0,
  input dut__core__ctrl___ctrlSignals_T_33_0,
  input dut__core__ctrl___ctrlSignals_T_45_0,
  input dut__core__ctrl___ctrlSignals_T_13_0,
  input dut__core__ctrl___ctrlSignals_T_53_0,
  input dut__core__ctrl___ctrlSignals_T_69_0,
  input dut__core__ctrl___ctrlSignals_T_3_0,
  input dut__core__ctrl___ctrlSignals_T_7_0,
  input dut__core__ctrl___ctrlSignals_T_73_0,
  input dut__core__ctrl___ctrlSignals_T_57_0,
  input dut__core__ctrl___ctrlSignals_T_61_0,
  input dut__icache___T_5_0,
  input dut__icache___wmask_T_0,
  input dut__icache___T_18_0,
  input dut__icache__io_cpu_req_valid_0,
  input dut__icache___T_25_0,
  input dut__icache___T_33_0,
  input dut__icache__wen_0,
  input dut__icache__is_alloc_reg_0,
  input dut__icache__read_wrap_out_0,
  input dut__icache___T_21_0,
  input dut__icache___T_11_0,
  input dut__icache___T_16_0,
  input dut__icache___T_0,
  input dut__icache__ren_0,
  input dut__icache___hit_T_2_0,
  input dut__icache___T_6_0,
  input dut__icache___io_nasti_ar_valid_T_0,
  input dut__icache___wen_T_0,
  input dut__icache__is_idle_0,
  input dut__icache___T_8_0,
  input dut__icache__is_write_0,
  input dut__icache___T_43_0,
  input dut__icache___T_20_0,
  input dut__icache___is_alloc_T_0,
  input dut__icache__read_count_0,
  input dut__icache___T_13_0,
  input dut__icache__io_cpu_resp_valid_0,
  input dut__icache___ren_T_0,
  input dut__icache___T_3_0,
  input dut__icache__ren_reg_0,
  input dut__icache___T_19_0,
  input dut__icache___T_51_0,
  input dut__icache___T_28_0,
  input dut__icache___T_9_0,
  input dut__icache___T_14_0,
  input dut__icache___T_4_0,
  input dut__icache___T_47_0,
  input dut__icache___T_15_0,
  input dut__icache___T_40_0,
  input dut__icache__is_alloc_0,
  input dut__icache__hit_0,
  input dut__icache___T_30_0,
  input dut__icache__is_read_0,
  input dut__icache___T_10_0,
  input dut__dcache___T_5_0,
  input dut__dcache___io_cpu_resp_valid_T_3_0,
  input dut__dcache___wmask_T_0,
  input dut__dcache___state_T_0,
  input dut__dcache__wen_0,
  input dut__dcache___T_33_0,
  input dut__dcache___T_44_0,
  input dut__dcache__read_wrap_out_0,
  input dut__dcache___T_21_0,
  input dut__dcache___T_16_0,
  input dut__dcache___ren_T_0,
  input dut__dcache__ren_0,
  input dut__dcache___hit_T_2_0,
  input dut__dcache___T_6_0,
  input dut__dcache___io_nasti_ar_valid_T_0,
  input dut__dcache___T_1_0,
  input dut__dcache___T_29_0,
  input dut__dcache__write_count_0,
  input dut__dcache___T_8_0,
  input dut__dcache__is_write_0,
  input dut__dcache___T_20_0,
  input dut__dcache___is_alloc_T_0,
  input dut__dcache__read_count_0,
  input dut__dcache__io_cpu_resp_valid_0,
  input dut__dcache___T_51_0,
  input dut__dcache___T_4_0,
  input dut__dcache___T_15_0,
  input dut__dcache___T_40_0,
  input dut__dcache__is_alloc_0,
  input dut__dcache__hit_0,
  input dut__dcache___T_30_0,
  input dut__dcache__is_read_0,
  input dut__dcache___T_35_0,
  input dut__dcache___T_10_0,
  input dut__dcache___T_18_0,
  input dut__dcache__io_cpu_req_valid_0,
  input dut__dcache___T_25_0,
  input dut__dcache__is_alloc_reg_0,
  input dut__dcache___T_11_0,
  input dut__dcache___T_0,
  input dut__dcache___io_cpu_resp_valid_T_2_0,
  input dut__dcache___wen_T_2_0,
  input dut__dcache__is_idle_0,
  input dut__dcache___T_43_0,
  input dut__dcache___T_13_0,
  input dut__dcache__write_wrap_out_0,
  input dut__dcache___T_3_0,
  input dut__dcache__ren_reg_0,
  input dut__dcache___T_19_0,
  input dut__dcache___T_28_0,
  input dut__dcache___T_9_0,
  input dut__dcache___T_14_0,
  input dut__dcache___T_47_0,
  input dut__arb___T_2_0,
  input dut__arb___T_13_0,
  input dut__arb___T_24_0,
  input dut__arb__io_dcache_ar_valid_0,
  input dut__arb___io_nasti_ar_valid_T_1_0,
  input dut__arb___T_20_0,
  input dut__arb___T_8_0,
  input dut__arb___io_dcache_b_valid_T_0,
  input dut__arb___T_5_0,
  input dut__arb___T_4_0,
  input dut__arb___io_icache_ar_ready_T_0,
  input dut__arb___T_10_0,
  input dut__arb___T_18_0,
  input dut__arb___io_nasti_aw_valid_T_0,
  input dut__arb___T_3_0,
  input dut__arb___io_icache_r_valid_T_0,
  input dut__arb___io_dcache_r_valid_T_0,
  input dut__arb___T_23_0,
  input dut__arb___io_nasti_w_valid_T_0
);
endmodule

