`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  wire [0:0] PI_clock = clock;
  reg [34:0] PI_io_inputs;
  Sodor5StageTop UUT (
    .clock(PI_clock),
    .io_inputs(PI_io_inputs)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$formal$Sodor5Stage_formal.\sv:453$1_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:454$2_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:455$3_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:456$4_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:457$5_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:458$6_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:459$7_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:460$8_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:461$9_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:462$10_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:463$11_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:464$12_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:465$13_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:466$14_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:467$15_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:468$16_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:469$17_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:470$18_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:471$19_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:472$20_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:473$21_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:474$22_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:475$23_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:476$24_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:477$25_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:478$26_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:479$27_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:480$28_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:481$29_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:482$30_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:483$31_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:484$32_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:485$33_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:486$34_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:487$35_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:488$36_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:489$37_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:490$38_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:491$39_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:492$40_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:493$41_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:494$42_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:495$43_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:496$44_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:497$45_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:498$46_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:499$47_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:500$48_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:501$49_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:502$50_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:503$51_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:504$52_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:505$53_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:506$54_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:507$55_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:508$56_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:509$57_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:510$58_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:511$59_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:512$60_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:513$61_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:514$62_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:515$63_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:516$64_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:517$65_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:518$66_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:519$67_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:520$68_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:521$69_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:522$70_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:523$71_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:524$72_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:525$73_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:526$74_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:527$75_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:528$76_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:529$77_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:530$78_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:531$79_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:532$80_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:533$81_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:534$82_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:535$83_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:536$84_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:537$85_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:538$86_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:539$87_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:540$88_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:541$89_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:542$90_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:543$91_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:544$92_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:545$93_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:546$94_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:547$95_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:548$96_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:549$97_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:550$98_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:551$99_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:552$100_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:553$101_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:554$102_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:555$103_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:556$104_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:557$105_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:558$106_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:559$107_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:560$108_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:561$109_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:562$110_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:563$111_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:564$112_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:565$113_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:566$114_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:567$115_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:568$116_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:569$117_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:570$118_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:571$119_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:572$120_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:573$121_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:574$122_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:575$123_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:576$124_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:577$125_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:578$126_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:579$127_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:580$128_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:581$129_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:582$130_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:583$131_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:584$132_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:585$133_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:586$134_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:587$135_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:588$136_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:589$137_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:590$138_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:591$139_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:592$140_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:593$141_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:594$142_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:595$143_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:596$144_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:597$145_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:598$146_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:599$147_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:600$148_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:601$149_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:602$150_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:603$151_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:604$152_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:605$153_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:606$154_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:607$155_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:608$156_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:609$157_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:610$158_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:611$159_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:612$160_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:613$161_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:614$162_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:615$163_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:616$164_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:617$165_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:618$166_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:619$167_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:620$168_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:621$169_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:622$170_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:623$171_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:624$172_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:625$173_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:626$174_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:627$175_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:628$176_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:629$177_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:630$178_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:631$179_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:632$180_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:633$181_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:634$182_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:635$183_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:636$184_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:637$185_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:638$186_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:639$187_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:640$188_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:641$189_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:642$190_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:643$191_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:644$192_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:645$193_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:646$194_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:647$195_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:648$196_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:649$197_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:650$198_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:651$199_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:652$200_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:653$201_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:654$202_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:655$203_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:656$204_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:657$205_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:658$206_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:659$207_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:660$208_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:661$209_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:662$210_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:663$211_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:664$212_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:665$213_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:666$214_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:667$215_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:668$216_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:669$217_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:670$218_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:671$219_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:672$220_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:673$221_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:674$222_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:675$223_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:676$224_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:677$225_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:678$226_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:679$227_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:680$228_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:681$229_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:682$230_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:683$231_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:684$232_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:685$233_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:686$234_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:687$235_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:688$236_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:689$237_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:690$238_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:691$239_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:692$240_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:693$241_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:694$242_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:695$243_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:696$244_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:697$245_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:698$246_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:699$247_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:700$248_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:701$249_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:702$250_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:703$251_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:704$252_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:705$253_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:706$254_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:707$255_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:708$256_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:709$257_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:710$258_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:711$259_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:712$260_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:713$261_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:714$262_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:715$263_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:716$264_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:717$265_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:718$266_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:719$267_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:720$268_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:721$269_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:722$270_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:723$271_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:724$272_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:725$273_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:726$274_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:727$275_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:728$276_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:729$277_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:730$278_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:731$279_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:732$280_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:733$281_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:734$282_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:735$283_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:736$284_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:737$285_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:738$286_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:739$287_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:740$288_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:741$289_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:742$290_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:743$291_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:744$292_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:745$293_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:746$294_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:747$295_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:748$296_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:749$297_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:750$298_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:751$299_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:752$300_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:753$301_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:754$302_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:755$303_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:756$304_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:757$305_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:758$306_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:759$307_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:760$308_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:761$309_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:762$310_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:763$311_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:764$312_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:765$313_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:766$314_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:767$315_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:768$316_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:769$317_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:770$318_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:771$319_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:772$320_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:773$321_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:774$322_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:775$323_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:776$324_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:777$325_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:778$326_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:779$327_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:780$328_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:781$329_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:782$330_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:783$331_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:784$332_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:785$333_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:786$334_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:787$335_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:788$336_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:789$337_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:790$338_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:791$339_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:792$340_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:793$341_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:794$342_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:795$343_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:796$344_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:797$345_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:798$346_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:799$347_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:800$348_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:801$349_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:802$350_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:803$351_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:804$352_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:805$353_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:806$354_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:807$355_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:808$356_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:809$357_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:810$358_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:811$359_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:812$360_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:813$361_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:814$362_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:815$363_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:816$364_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:817$365_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:818$366_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:819$367_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:820$368_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:821$369_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:822$370_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:823$371_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:824$372_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:825$373_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:826$374_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:827$375_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:828$376_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:829$377_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:830$378_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:831$379_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:832$380_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:833$381_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:834$382_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:835$383_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:836$384_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:837$385_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:838$386_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:839$387_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:840$388_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:841$389_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:842$390_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:843$391_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:844$392_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:845$393_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:846$394_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:847$395_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:848$396_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:849$397_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:850$398_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:851$399_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:852$400_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:853$401_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:854$402_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:855$403_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:856$404_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:857$405_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:858$406_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:859$407_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:860$408_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:861$409_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:862$410_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:863$411_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:864$412_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:865$413_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:866$414_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:867$415_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:868$416_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:869$417_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:870$418_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:871$419_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:872$420_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:873$421_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:874$422_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:875$423_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:876$424_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:877$425_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:878$426_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:879$427_CHECK  = 1'b0;
    // UUT.$formal$Sodor5Stage_formal.\sv:880$428_CHECK  = 1'b1;
    // UUT.$formal$Sodor5Stage_formal.\sv:888$429_EN  = 1'b0;
    UUT.bb.core.c._T_1152 = 1'b0;
    UUT.bb.core.c._T_1222 = 1'b0;
    UUT.bb.core.c._T_1225 = 1'b0;
    UUT.bb.core.c.exe_inst_is_load = 1'b1;
    UUT.bb.core.c.exe_reg_exception = 1'b0;
    UUT.bb.core.c.exe_reg_is_csr = 1'b0;
    UUT.bb.core.c.exe_reg_wbaddr = 5'b00001;
    UUT.bb.core.d.brjmp_offset = 32'b00000000000000000000000000000000;
    UUT.bb.core.d.csr._T_176 = 6'b010100;
    UUT.bb.core.d.csr._T_180 = 58'b0000000000000000000000000000000010000000000000010010001100;
    UUT.bb.core.d.csr._T_188 = 6'b111111;
    UUT.bb.core.d.csr._T_192 = 58'b0000000000000000000000000000000010000000000000010010001100;
    UUT.bb.core.d.csr._T_200 = 40'b0000000010000000000001000010001100000000;
    UUT.bb.core.d.csr._T_203 = 40'b0000000010000000000000000000000000000000;
    UUT.bb.core.d.csr._T_206 = 40'b0000000010000000000000010010001100010000;
    UUT.bb.core.d.csr._T_209 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_212 = 40'b0000000010000000000000100010010100000001;
    UUT.bb.core.d.csr._T_215 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_218 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_221 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_224 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_227 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_230 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_233 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_236 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_239 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_242 = 40'b0000000010000100000000000010001100000001;
    UUT.bb.core.d.csr._T_245 = 40'b0000000010000100000000000000010001000000;
    UUT.bb.core.d.csr._T_248 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_251 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_254 = 40'b0000000010000000000000010010010100000001;
    UUT.bb.core.d.csr._T_257 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_260 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_263 = 40'b0000000011000000000000000010001100000001;
    UUT.bb.core.d.csr._T_266 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_269 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_272 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_275 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_278 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_281 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_284 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_287 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_290 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr._T_293 = 40'b0000000010000000000000010010001100000001;
    UUT.bb.core.d.csr.reg_dcsr_ebreakm = 1'b1;
    UUT.bb.core.d.csr.reg_dcsr_step = 1'b0;
    UUT.bb.core.d.csr.reg_dpc = 32'b10000000000000010010001100000001;
    UUT.bb.core.d.csr.reg_dscratch = 32'b10000000000000010010001100000001;
    UUT.bb.core.d.csr.reg_mcause = 32'b10000000000000010010001100000001;
    UUT.bb.core.d.csr.reg_medeleg = 32'b10000000000010000000001100000001;
    UUT.bb.core.d.csr.reg_mepc = 32'b10000000000000010010001100000001;
    UUT.bb.core.d.csr.reg_mie_msip = 1'b0;
    UUT.bb.core.d.csr.reg_mie_mtip = 1'b1;
    UUT.bb.core.d.csr.reg_mip_msip = 1'b0;
    UUT.bb.core.d.csr.reg_mip_mtip = 1'b1;
    UUT.bb.core.d.csr.reg_mscratch = 32'b10000000000000010010001100000001;
    UUT.bb.core.d.csr.reg_mstatus_mie = 1'b0;
    UUT.bb.core.d.csr.reg_mstatus_mpie = 1'b0;
    UUT.bb.core.d.csr.reg_mtval = 32'b10000000000000010010001100000001;
    UUT.bb.core.d.dec_reg_inst = 32'b00000000000010010000000000000000;
    UUT.bb.core.d.dec_reg_pc = 32'b00000000000000000000000000000000;
    UUT.bb.core.d.exe_alu_op1 = 32'b00000000000000000000000000000000;
    UUT.bb.core.d.exe_reg_ctrl_alu_fun = 4'b0100;
    UUT.bb.core.d.exe_reg_ctrl_br_type = 4'b0000;
    UUT.bb.core.d.exe_reg_ctrl_csr_cmd = 3'b000;
    UUT.bb.core.d.exe_reg_ctrl_mem_fcn = 1'b0;
    UUT.bb.core.d.exe_reg_ctrl_mem_typ = 3'b000;
    UUT.bb.core.d.exe_reg_ctrl_mem_val = 1'b0;
    UUT.bb.core.d.exe_reg_ctrl_rf_wen = 1'b0;
    UUT.bb.core.d.exe_reg_ctrl_wb_sel = 2'b00;
    UUT.bb.core.d.exe_reg_inst = 32'b00000000000000000100000000110011;
    UUT.bb.core.d.exe_reg_pc = 32'b00000000000000000000000000000000;
    UUT.bb.core.d.exe_reg_rs2_data = 32'b00000000000000000000000000000001;
    UUT.bb.core.d.exe_reg_wbaddr = 5'b10010;
    UUT.bb.core.d.if_reg_pc = 32'b00000000000000000000000000000000;
    UUT.bb.core.d.mem_reg_alu_out = 32'b00000000000000000000000000000010;
    UUT.bb.core.d.mem_reg_ctrl_csr_cmd = 3'b000;
    UUT.bb.core.d.mem_reg_ctrl_mem_fcn = 1'b0;
    UUT.bb.core.d.mem_reg_ctrl_mem_typ = 3'b001;
    UUT.bb.core.d.mem_reg_ctrl_mem_val = 1'b0;
    UUT.bb.core.d.mem_reg_ctrl_rf_wen = 1'b1;
    UUT.bb.core.d.mem_reg_ctrl_wb_sel = 2'b11;
    UUT.bb.core.d.mem_reg_inst = 32'b11100000000000000000000000000000;
    UUT.bb.core.d.mem_reg_pc = 32'b00000000000000000000000000000000;
    UUT.bb.core.d.mem_reg_rs2_data = 32'b00000000000000000000000000000000;
    UUT.bb.core.d.mem_reg_wbaddr = 5'b00001;
    UUT.bb.core.d.regfile.mem_sparse.addresses_0_bits = 5'b00000;
    UUT.bb.core.d.regfile.mem_sparse.addresses_10_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_11_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_12_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_13_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_14_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_15_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_16_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_17_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_18_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_19_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_1_bits = 5'b00000;
    UUT.bb.core.d.regfile.mem_sparse.addresses_20_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_21_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_22_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_23_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_24_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_25_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_26_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_27_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_28_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_29_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_2_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_30_bits = 5'b10000;
    UUT.bb.core.d.regfile.mem_sparse.addresses_31_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_3_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_4_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_5_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_6_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_7_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_8_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.addresses_9_bits = 5'b00010;
    UUT.bb.core.d.regfile.mem_sparse.nextAddr = 6'b001000;
    UUT.bb.core.d.wb_reg_ctrl_rf_wen = 1'b1;
    UUT.bb.core.d.wb_reg_wbaddr = 5'b00001;
    UUT.bb.core.d.wb_reg_wbdata = 32'b00000000000000000000000000000000;
    UUT.bb.memory.async_data.mem_sparse.addresses_0_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse.addresses_10_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_11_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_12_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_13_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_14_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_15_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_16_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_17_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_18_bits = 21'b000000000000000001000;
    UUT.bb.memory.async_data.mem_sparse.addresses_19_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_1_bits = 21'b000000000000100100000;
    UUT.bb.memory.async_data.mem_sparse.addresses_20_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_21_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_22_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_23_bits = 21'b000000000000000000100;
    UUT.bb.memory.async_data.mem_sparse.addresses_24_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_25_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_26_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_27_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_28_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_29_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_2_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_30_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_31_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_3_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_4_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_5_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_6_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_7_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_8_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.addresses_9_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.nextAddr = 6'b010000;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_0_bits = 21'b010000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_10_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_11_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_12_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_13_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_14_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_15_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_16_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_17_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_18_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_19_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_1_bits = 21'b000000000000100000000;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_20_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_21_bits = 21'b000000000000000000100;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_22_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_23_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_24_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_25_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_26_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_27_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_28_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_29_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_2_bits = 21'b000000000000100100000;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_30_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_31_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_3_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_4_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_5_bits = 21'b000000000100000000000;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_6_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_7_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_8_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.addresses_9_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_0.nextAddr = 6'b000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_0_bits = 21'b000000001000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_10_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_11_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_12_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_13_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_14_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_15_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_16_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_17_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_18_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_19_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_1_bits = 21'b000000000000000000010;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_20_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_21_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_22_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_23_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_24_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_25_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_26_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_27_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_28_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_29_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_2_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_30_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_31_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_3_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_4_bits = 21'b000000000000100100000;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_5_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_6_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_7_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_8_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.addresses_9_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_1.nextAddr = 6'b010000;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_0_bits = 21'b000000000100000000010;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_10_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_11_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_12_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_13_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_14_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_15_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_16_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_17_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_18_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_19_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_1_bits = 21'b000000000000000000100;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_20_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_21_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_22_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_23_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_24_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_25_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_26_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_27_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_28_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_29_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_2_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_30_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_31_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_3_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_4_bits = 21'b000000100000000000000;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_5_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_6_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_7_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_8_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.addresses_9_bits = 21'b000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse_2.nextAddr = 6'b001000;
    UUT.is_meta_reset_phase = 1'b1;
    UUT.is_reset_phase = 1'b0;
    UUT.bb.core.d.regfile.mem_sparse.mem[5'b00001] = 32'b10000000000000000000000000000000;
    UUT.bb.core.d.regfile.mem_sparse.mem[5'b00000] = 32'b00000000000000000000000000000000;
    UUT.bb.core.d.regfile.mem_sparse.mem[5'b11111] = 32'b00000000000000000000000000000001;
    UUT.bb.memory.async_data.mem_sparse.mem[5'b00000] = 8'b01000110;
    UUT.bb.memory.async_data.mem_sparse.mem[5'b11111] = 8'b00000001;
    UUT.bb.memory.async_data.mem_sparse_0.mem[5'b00000] = 8'b00000000;
    UUT.bb.memory.async_data.mem_sparse_0.mem[5'b11111] = 8'b00000001;
    UUT.bb.memory.async_data.mem_sparse_1.mem[5'b00001] = 8'b00000100;
    UUT.bb.memory.async_data.mem_sparse_1.mem[5'b11111] = 8'b00000001;
    UUT.bb.memory.async_data.mem_sparse_1.mem[5'b00000] = 8'b00000000;
    UUT.bb.memory.async_data.mem_sparse_2.mem[5'b00000] = 8'b00000000;
    UUT.bb.memory.async_data.mem_sparse_2.mem[5'b11111] = 8'b00000000;

    // state 0
    PI_io_inputs = 35'b00000000000000000000000000000000000;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_io_inputs <= 35'b00000000000000000000000000000000010;
    end

    // state 2
    if (cycle == 1) begin
      PI_io_inputs <= 35'b00000100010001000000001000010111010;
    end

    // state 3
    if (cycle == 2) begin
      PI_io_inputs <= 35'b00000000010000100001001000000011010;
    end

    // state 4
    if (cycle == 3) begin
      PI_io_inputs <= 35'b10000000000000000000000000000010010;
    end

    // state 5
    if (cycle == 4) begin
      PI_io_inputs <= 35'b00000000000000000000000000000000000;
    end

    genclock <= cycle < 5;
    cycle <= cycle + 1;
  end
endmodule
