`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  reg [34:0] PI_io_inputs;
  wire [0:0] PI_clock = clock;
  Sodor3StageTop UUT (
    .io_inputs(PI_io_inputs),
    .clock(PI_clock)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$formal$Sodor3Stage_formal.\sv:399$1_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:400$2_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:401$3_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:402$4_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:403$5_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:404$6_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:405$7_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:406$8_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:407$9_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:408$10_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:409$11_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:410$12_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:411$13_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:412$14_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:413$15_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:414$16_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:415$17_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:416$18_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:417$19_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:418$20_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:419$21_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:420$22_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:421$23_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:422$24_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:423$25_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:424$26_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:425$27_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:426$28_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:427$29_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:428$30_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:429$31_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:430$32_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:431$33_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:432$34_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:433$35_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:434$36_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:435$37_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:436$38_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:437$39_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:438$40_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:439$41_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:440$42_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:441$43_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:442$44_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:443$45_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:444$46_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:445$47_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:446$48_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:447$49_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:448$50_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:449$51_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:450$52_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:451$53_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:452$54_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:453$55_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:454$56_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:455$57_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:456$58_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:457$59_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:458$60_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:459$61_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:460$62_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:461$63_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:462$64_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:463$65_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:464$66_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:465$67_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:466$68_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:467$69_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:468$70_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:469$71_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:470$72_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:471$73_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:472$74_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:473$75_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:474$76_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:475$77_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:476$78_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:477$79_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:478$80_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:479$81_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:480$82_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:481$83_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:482$84_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:483$85_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:484$86_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:485$87_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:486$88_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:487$89_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:488$90_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:489$91_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:490$92_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:491$93_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:492$94_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:493$95_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:494$96_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:495$97_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:496$98_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:497$99_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:498$100_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:499$101_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:500$102_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:501$103_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:502$104_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:503$105_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:504$106_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:505$107_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:506$108_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:507$109_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:508$110_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:509$111_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:510$112_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:511$113_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:512$114_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:513$115_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:514$116_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:515$117_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:516$118_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:517$119_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:518$120_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:519$121_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:520$122_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:521$123_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:522$124_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:523$125_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:524$126_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:525$127_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:526$128_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:527$129_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:528$130_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:529$131_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:530$132_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:531$133_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:532$134_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:533$135_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:534$136_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:535$137_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:536$138_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:537$139_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:538$140_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:539$141_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:540$142_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:541$143_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:542$144_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:543$145_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:544$146_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:545$147_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:546$148_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:547$149_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:548$150_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:549$151_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:550$152_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:551$153_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:552$154_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:553$155_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:554$156_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:555$157_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:556$158_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:557$159_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:558$160_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:559$161_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:560$162_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:561$163_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:562$164_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:563$165_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:564$166_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:565$167_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:566$168_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:567$169_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:568$170_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:569$171_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:570$172_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:571$173_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:572$174_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:573$175_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:574$176_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:575$177_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:576$178_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:577$179_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:578$180_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:579$181_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:580$182_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:581$183_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:582$184_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:583$185_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:584$186_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:585$187_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:586$188_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:587$189_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:588$190_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:589$191_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:590$192_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:591$193_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:592$194_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:593$195_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:594$196_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:595$197_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:596$198_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:597$199_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:598$200_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:599$201_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:600$202_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:601$203_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:602$204_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:603$205_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:604$206_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:605$207_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:606$208_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:607$209_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:608$210_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:609$211_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:610$212_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:611$213_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:612$214_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:613$215_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:614$216_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:615$217_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:616$218_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:617$219_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:618$220_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:619$221_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:620$222_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:621$223_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:622$224_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:623$225_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:624$226_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:625$227_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:626$228_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:627$229_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:628$230_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:629$231_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:630$232_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:631$233_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:632$234_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:633$235_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:634$236_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:635$237_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:636$238_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:637$239_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:638$240_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:639$241_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:640$242_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:641$243_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:642$244_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:643$245_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:644$246_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:645$247_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:646$248_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:647$249_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:648$250_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:649$251_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:650$252_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:651$253_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:652$254_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:653$255_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:654$256_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:655$257_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:656$258_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:657$259_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:658$260_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:659$261_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:660$262_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:661$263_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:662$264_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:663$265_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:664$266_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:665$267_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:666$268_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:667$269_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:668$270_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:669$271_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:670$272_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:671$273_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:672$274_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:673$275_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:674$276_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:675$277_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:676$278_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:677$279_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:678$280_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:679$281_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:680$282_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:681$283_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:682$284_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:683$285_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:684$286_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:685$287_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:686$288_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:687$289_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:688$290_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:689$291_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:690$292_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:691$293_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:692$294_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:693$295_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:694$296_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:695$297_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:696$298_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:697$299_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:698$300_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:699$301_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:700$302_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:701$303_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:702$304_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:703$305_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:704$306_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:705$307_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:706$308_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:707$309_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:708$310_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:709$311_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:710$312_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:711$313_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:712$314_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:713$315_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:714$316_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:715$317_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:716$318_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:717$319_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:718$320_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:719$321_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:720$322_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:721$323_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:722$324_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:723$325_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:724$326_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:725$327_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:726$328_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:727$329_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:728$330_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:729$331_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:730$332_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:731$333_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:732$334_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:733$335_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:734$336_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:735$337_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:736$338_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:737$339_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:738$340_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:739$341_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:740$342_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:741$343_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:742$344_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:743$345_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:744$346_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:745$347_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:746$348_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:747$349_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:748$350_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:749$351_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:750$352_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:751$353_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:752$354_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:753$355_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:754$356_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:755$357_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:756$358_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:757$359_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:758$360_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:759$361_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:760$362_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:761$363_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:762$364_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:763$365_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:764$366_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:765$367_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:766$368_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:767$369_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:768$370_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:769$371_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:770$372_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:771$373_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:772$374_CHECK  = 1'b0;
    // UUT.$formal$Sodor3Stage_formal.\sv:780$375_EN  = 1'b0;
    UUT.bb.core.cpath._T_1028 = 1'b0;
    UUT.bb.core.dpath._T_246 = 1'b0;
    UUT.bb.core.dpath.csr._T_176 = 6'b000000;
    UUT.bb.core.dpath.csr._T_180 = 58'b0000000000000000000000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_188 = 6'b000000;
    UUT.bb.core.dpath.csr._T_192 = 58'b0000000000000000000000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_200 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_203 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_206 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_209 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_212 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_215 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_218 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_221 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_224 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_227 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_230 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_233 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_236 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_239 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_242 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_245 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_248 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_251 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_254 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_257 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_260 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_263 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_266 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_269 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_272 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_275 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_278 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_281 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_284 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_287 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_290 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr._T_293 = 40'b0000000000000000000000000000000000000000;
    UUT.bb.core.dpath.csr.reg_dcsr_ebreakm = 1'b0;
    UUT.bb.core.dpath.csr.reg_dcsr_step = 1'b0;
    UUT.bb.core.dpath.csr.reg_dpc = 32'b00000000000000000000000000000000;
    UUT.bb.core.dpath.csr.reg_dscratch = 32'b00000000000000000000000000000000;
    UUT.bb.core.dpath.csr.reg_mcause = 32'b00000000000000000000000000000000;
    UUT.bb.core.dpath.csr.reg_medeleg = 32'b00000000000000000000000000000000;
    UUT.bb.core.dpath.csr.reg_mepc = 32'b00000000000000000000000000000000;
    UUT.bb.core.dpath.csr.reg_mie_msip = 1'b0;
    UUT.bb.core.dpath.csr.reg_mie_mtip = 1'b0;
    UUT.bb.core.dpath.csr.reg_mip_msip = 1'b0;
    UUT.bb.core.dpath.csr.reg_mip_mtip = 1'b0;
    UUT.bb.core.dpath.csr.reg_mscratch = 32'b00000000000000000000000000000000;
    UUT.bb.core.dpath.csr.reg_mstatus_mie = 1'b0;
    UUT.bb.core.dpath.csr.reg_mstatus_mpie = 1'b0;
    UUT.bb.core.dpath.csr.reg_mtval = 32'b00000000000000000000000000000000;
    UUT.bb.core.dpath.mem_sparse.addresses_0_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_0_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_10_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_10_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_11_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_11_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_12_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_12_valid = 1'b1;
    UUT.bb.core.dpath.mem_sparse.addresses_13_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_13_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_14_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_14_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_15_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_15_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_16_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_16_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_17_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_17_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_18_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_18_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_19_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_19_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_1_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_1_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_20_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_20_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_21_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_21_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_22_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_22_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_23_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_23_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_24_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_24_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_25_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_25_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_26_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_26_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_27_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_27_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_28_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_28_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_29_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_29_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_2_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_2_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_30_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_30_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_31_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_31_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_3_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_3_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_4_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_4_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_5_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_5_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_6_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_6_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_7_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_7_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_8_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_8_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.addresses_9_bits = 5'b10001;
    UUT.bb.core.dpath.mem_sparse.addresses_9_valid = 1'b0;
    UUT.bb.core.dpath.mem_sparse.nextAddr = 6'b000000;
    UUT.bb.core.dpath.wb_reg_alu = 32'b00000000000000001111111111111111;
    UUT.bb.core.dpath.wb_reg_csr_addr = 12'b000000000000;
    UUT.bb.core.dpath.wb_reg_ctrl_bypassable = 1'b1;
    UUT.bb.core.dpath.wb_reg_ctrl_csr_cmd = 3'b000;
    UUT.bb.core.dpath.wb_reg_ctrl_rf_wen = 1'b1;
    UUT.bb.core.dpath.wb_reg_ctrl_wb_sel = 2'b00;
    UUT.bb.core.dpath.wb_reg_valid = 1'b0;
    UUT.bb.core.dpath.wb_reg_wbaddr = 5'b10000;
    UUT.bb.core.frontend.exe_reg_inst = 32'b00000001000010001000111000100011;
    UUT.bb.core.frontend.exe_reg_pc = 32'b11111111111111111111111111111111;
    UUT.bb.core.frontend.exe_reg_valid = 1'b1;
    UUT.bb.core.frontend.if_reg_pc = 32'b00000000000000000000000000000000;
    UUT.bb.core.frontend.if_reg_valid = 1'b0;
    UUT.bb.memory.req_typi = 3'b000;
    UUT.bb.memory.sync_data.mem_sparse.addresses_0_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_10_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_11_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_12_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_13_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_14_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_15_bits = 21'b111111111111111111111;
    UUT.bb.memory.sync_data.mem_sparse.addresses_16_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_17_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_18_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_19_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_1_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_20_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_21_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_22_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_23_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_24_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_25_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_26_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_27_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_28_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_29_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_2_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_30_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_31_bits = 21'b111111111111111111111;
    UUT.bb.memory.sync_data.mem_sparse.addresses_3_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_4_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_5_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_6_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_7_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_8_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.addresses_9_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse.nextAddr = 6'b111111;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_0_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_10_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_11_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_12_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_13_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_14_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_15_bits = 21'b111111111111111111111;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_16_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_17_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_18_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_19_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_1_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_20_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_21_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_22_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_23_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_24_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_25_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_26_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_27_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_28_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_29_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_2_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_30_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_31_bits = 21'b111111111111111111111;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_3_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_4_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_5_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_6_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_7_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_8_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.addresses_9_bits = 21'b111111111111111111110;
    UUT.bb.memory.sync_data.mem_sparse_0.nextAddr = 6'b111111;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_0_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_10_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_11_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_12_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_13_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_14_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_15_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_16_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_17_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_18_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_19_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_1_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_20_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_21_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_22_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_23_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_24_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_25_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_26_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_27_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_28_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_29_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_2_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_30_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_31_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_3_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_4_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_5_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_6_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_7_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_8_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.addresses_9_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_1.nextAddr = 6'b000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_0_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_10_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_11_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_12_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_13_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_14_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_15_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_16_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_17_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_18_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_19_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_1_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_20_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_21_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_22_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_23_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_24_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_25_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_26_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_27_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_28_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_29_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_2_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_30_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_31_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_3_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_4_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_5_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_6_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_7_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_8_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.addresses_9_bits = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.mem_sparse_2.nextAddr = 6'b000000;
    UUT.bb.memory.sync_data.underlying_0__T_54_addr_pipe_0 = 21'b111111111111111111111;
    UUT.bb.memory.sync_data.underlying_1__T_54_addr_pipe_0 = 21'b111111111111111111111;
    UUT.bb.memory.sync_data.underlying_2__T_54_addr_pipe_0 = 21'b000000000000000000000;
    UUT.bb.memory.sync_data.underlying_3__T_54_addr_pipe_0 = 21'b000000000000000000000;
    UUT.is_meta_reset_phase = 1'b1;
    UUT.is_reset_phase = 1'b0;
    UUT.bb.core.dpath.mem_sparse.mem[5'b00000] = 32'b11111111111111111111111111111111;
    UUT.bb.core.dpath.mem_sparse.mem[5'b01100] = 32'b11111111111111111111111111100000;
    UUT.bb.memory.sync_data.mem_sparse.mem[5'b11111] = 8'b11111111;
    UUT.bb.memory.sync_data.mem_sparse_0.mem[5'b11111] = 8'b11111111;
    UUT.bb.memory.sync_data.mem_sparse_1.mem[5'b11111] = 8'b00000000;
    UUT.bb.memory.sync_data.mem_sparse_2.mem[5'b11111] = 8'b00000000;

    // state 0
    PI_io_inputs = 35'b00000000000000000000000000000000000;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_io_inputs <= 35'b10111001111000000101000001110011000;
    end

    // state 2
    if (cycle == 1) begin
      PI_io_inputs <= 35'b00000000000000000000000001100111000;
    end

    // state 3
    if (cycle == 2) begin
      PI_io_inputs <= 35'b00000001111111111101111111110011000;
    end

    // state 4
    if (cycle == 3) begin
      PI_io_inputs <= 35'b00000000000000000000000000000000000;
    end

    genclock <= cycle < 4;
    cycle <= cycle + 1;
  end
endmodule
